magic
tech sky130A
magscale 1 2
timestamp 1712816020
<< pwell >>
rect -686 -300 686 300
<< nmos >>
rect -500 -100 500 100
<< ndiff >>
rect -558 85 -500 100
rect -558 51 -546 85
rect -512 51 -500 85
rect -558 17 -500 51
rect -558 -17 -546 17
rect -512 -17 -500 17
rect -558 -51 -500 -17
rect -558 -85 -546 -51
rect -512 -85 -500 -51
rect -558 -100 -500 -85
rect 500 85 558 100
rect 500 51 512 85
rect 546 51 558 85
rect 500 17 558 51
rect 500 -17 512 17
rect 546 -17 558 17
rect 500 -51 558 -17
rect 500 -85 512 -51
rect 546 -85 558 -51
rect 500 -100 558 -85
<< ndiffc >>
rect -546 51 -512 85
rect -546 -17 -512 17
rect -546 -85 -512 -51
rect 512 51 546 85
rect 512 -17 546 17
rect 512 -85 546 -51
<< psubdiff >>
rect -660 240 -561 274
rect -527 240 -493 274
rect -459 240 -425 274
rect -391 240 -357 274
rect -323 240 -289 274
rect -255 240 -221 274
rect -187 240 -153 274
rect -119 240 -85 274
rect -51 240 -17 274
rect 17 240 51 274
rect 85 240 119 274
rect 153 240 187 274
rect 221 240 255 274
rect 289 240 323 274
rect 357 240 391 274
rect 425 240 459 274
rect 493 240 527 274
rect 561 240 660 274
rect -660 153 -626 240
rect -660 85 -626 119
rect 626 153 660 240
rect -660 17 -626 51
rect -660 -51 -626 -17
rect -660 -119 -626 -85
rect 626 85 660 119
rect 626 17 660 51
rect 626 -51 660 -17
rect -660 -240 -626 -153
rect 626 -119 660 -85
rect 626 -240 660 -153
rect -660 -274 -561 -240
rect -527 -274 -493 -240
rect -459 -274 -425 -240
rect -391 -274 -357 -240
rect -323 -274 -289 -240
rect -255 -274 -221 -240
rect -187 -274 -153 -240
rect -119 -274 -85 -240
rect -51 -274 -17 -240
rect 17 -274 51 -240
rect 85 -274 119 -240
rect 153 -274 187 -240
rect 221 -274 255 -240
rect 289 -274 323 -240
rect 357 -274 391 -240
rect 425 -274 459 -240
rect 493 -274 527 -240
rect 561 -274 660 -240
<< psubdiffcont >>
rect -561 240 -527 274
rect -493 240 -459 274
rect -425 240 -391 274
rect -357 240 -323 274
rect -289 240 -255 274
rect -221 240 -187 274
rect -153 240 -119 274
rect -85 240 -51 274
rect -17 240 17 274
rect 51 240 85 274
rect 119 240 153 274
rect 187 240 221 274
rect 255 240 289 274
rect 323 240 357 274
rect 391 240 425 274
rect 459 240 493 274
rect 527 240 561 274
rect -660 119 -626 153
rect 626 119 660 153
rect -660 51 -626 85
rect -660 -17 -626 17
rect -660 -85 -626 -51
rect 626 51 660 85
rect 626 -17 660 17
rect 626 -85 660 -51
rect -660 -153 -626 -119
rect 626 -153 660 -119
rect -561 -274 -527 -240
rect -493 -274 -459 -240
rect -425 -274 -391 -240
rect -357 -274 -323 -240
rect -289 -274 -255 -240
rect -221 -274 -187 -240
rect -153 -274 -119 -240
rect -85 -274 -51 -240
rect -17 -274 17 -240
rect 51 -274 85 -240
rect 119 -274 153 -240
rect 187 -274 221 -240
rect 255 -274 289 -240
rect 323 -274 357 -240
rect 391 -274 425 -240
rect 459 -274 493 -240
rect 527 -274 561 -240
<< poly >>
rect -500 172 500 188
rect -500 138 -459 172
rect -425 138 -391 172
rect -357 138 -323 172
rect -289 138 -255 172
rect -221 138 -187 172
rect -153 138 -119 172
rect -85 138 -51 172
rect -17 138 17 172
rect 51 138 85 172
rect 119 138 153 172
rect 187 138 221 172
rect 255 138 289 172
rect 323 138 357 172
rect 391 138 425 172
rect 459 138 500 172
rect -500 100 500 138
rect -500 -138 500 -100
rect -500 -172 -459 -138
rect -425 -172 -391 -138
rect -357 -172 -323 -138
rect -289 -172 -255 -138
rect -221 -172 -187 -138
rect -153 -172 -119 -138
rect -85 -172 -51 -138
rect -17 -172 17 -138
rect 51 -172 85 -138
rect 119 -172 153 -138
rect 187 -172 221 -138
rect 255 -172 289 -138
rect 323 -172 357 -138
rect 391 -172 425 -138
rect 459 -172 500 -138
rect -500 -188 500 -172
<< polycont >>
rect -459 138 -425 172
rect -391 138 -357 172
rect -323 138 -289 172
rect -255 138 -221 172
rect -187 138 -153 172
rect -119 138 -85 172
rect -51 138 -17 172
rect 17 138 51 172
rect 85 138 119 172
rect 153 138 187 172
rect 221 138 255 172
rect 289 138 323 172
rect 357 138 391 172
rect 425 138 459 172
rect -459 -172 -425 -138
rect -391 -172 -357 -138
rect -323 -172 -289 -138
rect -255 -172 -221 -138
rect -187 -172 -153 -138
rect -119 -172 -85 -138
rect -51 -172 -17 -138
rect 17 -172 51 -138
rect 85 -172 119 -138
rect 153 -172 187 -138
rect 221 -172 255 -138
rect 289 -172 323 -138
rect 357 -172 391 -138
rect 425 -172 459 -138
<< locali >>
rect -660 240 -561 274
rect -527 240 -493 274
rect -459 240 -425 274
rect -391 240 -357 274
rect -323 240 -289 274
rect -255 240 -221 274
rect -187 240 -153 274
rect -119 240 -85 274
rect -51 240 -17 274
rect 17 240 51 274
rect 85 240 119 274
rect 153 240 187 274
rect 221 240 255 274
rect 289 240 323 274
rect 357 240 391 274
rect 425 240 459 274
rect 493 240 527 274
rect 561 240 660 274
rect -660 153 -626 240
rect -500 138 -459 172
rect -415 138 -391 172
rect -343 138 -323 172
rect -271 138 -255 172
rect -199 138 -187 172
rect -127 138 -119 172
rect -55 138 -51 172
rect 51 138 55 172
rect 119 138 127 172
rect 187 138 199 172
rect 255 138 271 172
rect 323 138 343 172
rect 391 138 415 172
rect 459 138 500 172
rect 626 153 660 240
rect -660 85 -626 119
rect -660 17 -626 51
rect -660 -51 -626 -17
rect -660 -119 -626 -85
rect -546 85 -512 104
rect -546 17 -512 19
rect -546 -19 -512 -17
rect -546 -104 -512 -85
rect 512 85 546 104
rect 512 17 546 19
rect 512 -19 546 -17
rect 512 -104 546 -85
rect 626 85 660 119
rect 626 17 660 51
rect 626 -51 660 -17
rect 626 -119 660 -85
rect -660 -240 -626 -153
rect -500 -172 -459 -138
rect -415 -172 -391 -138
rect -343 -172 -323 -138
rect -271 -172 -255 -138
rect -199 -172 -187 -138
rect -127 -172 -119 -138
rect -55 -172 -51 -138
rect 51 -172 55 -138
rect 119 -172 127 -138
rect 187 -172 199 -138
rect 255 -172 271 -138
rect 323 -172 343 -138
rect 391 -172 415 -138
rect 459 -172 500 -138
rect 626 -240 660 -153
rect -660 -274 -561 -240
rect -527 -274 -493 -240
rect -459 -274 -425 -240
rect -391 -274 -357 -240
rect -323 -274 -289 -240
rect -255 -274 -221 -240
rect -187 -274 -153 -240
rect -119 -274 -85 -240
rect -51 -274 -17 -240
rect 17 -274 51 -240
rect 85 -274 119 -240
rect 153 -274 187 -240
rect 221 -274 255 -240
rect 289 -274 323 -240
rect 357 -274 391 -240
rect 425 -274 459 -240
rect 493 -274 527 -240
rect 561 -274 660 -240
<< viali >>
rect -449 138 -425 172
rect -425 138 -415 172
rect -377 138 -357 172
rect -357 138 -343 172
rect -305 138 -289 172
rect -289 138 -271 172
rect -233 138 -221 172
rect -221 138 -199 172
rect -161 138 -153 172
rect -153 138 -127 172
rect -89 138 -85 172
rect -85 138 -55 172
rect -17 138 17 172
rect 55 138 85 172
rect 85 138 89 172
rect 127 138 153 172
rect 153 138 161 172
rect 199 138 221 172
rect 221 138 233 172
rect 271 138 289 172
rect 289 138 305 172
rect 343 138 357 172
rect 357 138 377 172
rect 415 138 425 172
rect 425 138 449 172
rect -546 51 -512 53
rect -546 19 -512 51
rect -546 -51 -512 -19
rect -546 -53 -512 -51
rect 512 51 546 53
rect 512 19 546 51
rect 512 -51 546 -19
rect 512 -53 546 -51
rect -449 -172 -425 -138
rect -425 -172 -415 -138
rect -377 -172 -357 -138
rect -357 -172 -343 -138
rect -305 -172 -289 -138
rect -289 -172 -271 -138
rect -233 -172 -221 -138
rect -221 -172 -199 -138
rect -161 -172 -153 -138
rect -153 -172 -127 -138
rect -89 -172 -85 -138
rect -85 -172 -55 -138
rect -17 -172 17 -138
rect 55 -172 85 -138
rect 85 -172 89 -138
rect 127 -172 153 -138
rect 153 -172 161 -138
rect 199 -172 221 -138
rect 221 -172 233 -138
rect 271 -172 289 -138
rect 289 -172 305 -138
rect 343 -172 357 -138
rect 357 -172 377 -138
rect 415 -172 425 -138
rect 425 -172 449 -138
<< metal1 >>
rect -496 172 496 178
rect -496 138 -449 172
rect -415 138 -377 172
rect -343 138 -305 172
rect -271 138 -233 172
rect -199 138 -161 172
rect -127 138 -89 172
rect -55 138 -17 172
rect 17 138 55 172
rect 89 138 127 172
rect 161 138 199 172
rect 233 138 271 172
rect 305 138 343 172
rect 377 138 415 172
rect 449 138 496 172
rect -496 132 496 138
rect -552 53 -506 100
rect -552 19 -546 53
rect -512 19 -506 53
rect -552 -19 -506 19
rect -552 -53 -546 -19
rect -512 -53 -506 -19
rect -552 -100 -506 -53
rect 506 53 552 100
rect 506 19 512 53
rect 546 19 552 53
rect 506 -19 552 19
rect 506 -53 512 -19
rect 546 -53 552 -19
rect 506 -100 552 -53
rect -496 -138 496 -132
rect -496 -172 -449 -138
rect -415 -172 -377 -138
rect -343 -172 -305 -138
rect -271 -172 -233 -138
rect -199 -172 -161 -138
rect -127 -172 -89 -138
rect -55 -172 -17 -138
rect 17 -172 55 -138
rect 89 -172 127 -138
rect 161 -172 199 -138
rect 233 -172 271 -138
rect 305 -172 343 -138
rect 377 -172 415 -138
rect 449 -172 496 -138
rect -496 -178 496 -172
<< properties >>
string FIXED_BBOX -642 -256 642 256
<< end >>
