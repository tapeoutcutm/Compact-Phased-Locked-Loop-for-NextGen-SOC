magic
tech sky130A
magscale 1 2
timestamp 1712816020
<< error_p >>
rect -29 681 29 687
rect -29 647 -17 681
rect -29 641 29 647
rect -29 -647 29 -641
rect -29 -681 -17 -647
rect -29 -687 29 -681
<< nwell >>
rect -226 -819 226 819
<< pmos >>
rect -30 -600 30 600
<< pdiff >>
rect -88 561 -30 600
rect -88 527 -76 561
rect -42 527 -30 561
rect -88 493 -30 527
rect -88 459 -76 493
rect -42 459 -30 493
rect -88 425 -30 459
rect -88 391 -76 425
rect -42 391 -30 425
rect -88 357 -30 391
rect -88 323 -76 357
rect -42 323 -30 357
rect -88 289 -30 323
rect -88 255 -76 289
rect -42 255 -30 289
rect -88 221 -30 255
rect -88 187 -76 221
rect -42 187 -30 221
rect -88 153 -30 187
rect -88 119 -76 153
rect -42 119 -30 153
rect -88 85 -30 119
rect -88 51 -76 85
rect -42 51 -30 85
rect -88 17 -30 51
rect -88 -17 -76 17
rect -42 -17 -30 17
rect -88 -51 -30 -17
rect -88 -85 -76 -51
rect -42 -85 -30 -51
rect -88 -119 -30 -85
rect -88 -153 -76 -119
rect -42 -153 -30 -119
rect -88 -187 -30 -153
rect -88 -221 -76 -187
rect -42 -221 -30 -187
rect -88 -255 -30 -221
rect -88 -289 -76 -255
rect -42 -289 -30 -255
rect -88 -323 -30 -289
rect -88 -357 -76 -323
rect -42 -357 -30 -323
rect -88 -391 -30 -357
rect -88 -425 -76 -391
rect -42 -425 -30 -391
rect -88 -459 -30 -425
rect -88 -493 -76 -459
rect -42 -493 -30 -459
rect -88 -527 -30 -493
rect -88 -561 -76 -527
rect -42 -561 -30 -527
rect -88 -600 -30 -561
rect 30 561 88 600
rect 30 527 42 561
rect 76 527 88 561
rect 30 493 88 527
rect 30 459 42 493
rect 76 459 88 493
rect 30 425 88 459
rect 30 391 42 425
rect 76 391 88 425
rect 30 357 88 391
rect 30 323 42 357
rect 76 323 88 357
rect 30 289 88 323
rect 30 255 42 289
rect 76 255 88 289
rect 30 221 88 255
rect 30 187 42 221
rect 76 187 88 221
rect 30 153 88 187
rect 30 119 42 153
rect 76 119 88 153
rect 30 85 88 119
rect 30 51 42 85
rect 76 51 88 85
rect 30 17 88 51
rect 30 -17 42 17
rect 76 -17 88 17
rect 30 -51 88 -17
rect 30 -85 42 -51
rect 76 -85 88 -51
rect 30 -119 88 -85
rect 30 -153 42 -119
rect 76 -153 88 -119
rect 30 -187 88 -153
rect 30 -221 42 -187
rect 76 -221 88 -187
rect 30 -255 88 -221
rect 30 -289 42 -255
rect 76 -289 88 -255
rect 30 -323 88 -289
rect 30 -357 42 -323
rect 76 -357 88 -323
rect 30 -391 88 -357
rect 30 -425 42 -391
rect 76 -425 88 -391
rect 30 -459 88 -425
rect 30 -493 42 -459
rect 76 -493 88 -459
rect 30 -527 88 -493
rect 30 -561 42 -527
rect 76 -561 88 -527
rect 30 -600 88 -561
<< pdiffc >>
rect -76 527 -42 561
rect -76 459 -42 493
rect -76 391 -42 425
rect -76 323 -42 357
rect -76 255 -42 289
rect -76 187 -42 221
rect -76 119 -42 153
rect -76 51 -42 85
rect -76 -17 -42 17
rect -76 -85 -42 -51
rect -76 -153 -42 -119
rect -76 -221 -42 -187
rect -76 -289 -42 -255
rect -76 -357 -42 -323
rect -76 -425 -42 -391
rect -76 -493 -42 -459
rect -76 -561 -42 -527
rect 42 527 76 561
rect 42 459 76 493
rect 42 391 76 425
rect 42 323 76 357
rect 42 255 76 289
rect 42 187 76 221
rect 42 119 76 153
rect 42 51 76 85
rect 42 -17 76 17
rect 42 -85 76 -51
rect 42 -153 76 -119
rect 42 -221 76 -187
rect 42 -289 76 -255
rect 42 -357 76 -323
rect 42 -425 76 -391
rect 42 -493 76 -459
rect 42 -561 76 -527
<< nsubdiff >>
rect -190 749 -85 783
rect -51 749 -17 783
rect 17 749 51 783
rect 85 749 190 783
rect -190 663 -156 749
rect 156 663 190 749
rect -190 595 -156 629
rect -190 527 -156 561
rect -190 459 -156 493
rect -190 391 -156 425
rect -190 323 -156 357
rect -190 255 -156 289
rect -190 187 -156 221
rect -190 119 -156 153
rect -190 51 -156 85
rect -190 -17 -156 17
rect -190 -85 -156 -51
rect -190 -153 -156 -119
rect -190 -221 -156 -187
rect -190 -289 -156 -255
rect -190 -357 -156 -323
rect -190 -425 -156 -391
rect -190 -493 -156 -459
rect -190 -561 -156 -527
rect -190 -629 -156 -595
rect 156 595 190 629
rect 156 527 190 561
rect 156 459 190 493
rect 156 391 190 425
rect 156 323 190 357
rect 156 255 190 289
rect 156 187 190 221
rect 156 119 190 153
rect 156 51 190 85
rect 156 -17 190 17
rect 156 -85 190 -51
rect 156 -153 190 -119
rect 156 -221 190 -187
rect 156 -289 190 -255
rect 156 -357 190 -323
rect 156 -425 190 -391
rect 156 -493 190 -459
rect 156 -561 190 -527
rect 156 -629 190 -595
rect -190 -749 -156 -663
rect 156 -749 190 -663
rect -190 -783 -85 -749
rect -51 -783 -17 -749
rect 17 -783 51 -749
rect 85 -783 190 -749
<< nsubdiffcont >>
rect -85 749 -51 783
rect -17 749 17 783
rect 51 749 85 783
rect -190 629 -156 663
rect 156 629 190 663
rect -190 561 -156 595
rect -190 493 -156 527
rect -190 425 -156 459
rect -190 357 -156 391
rect -190 289 -156 323
rect -190 221 -156 255
rect -190 153 -156 187
rect -190 85 -156 119
rect -190 17 -156 51
rect -190 -51 -156 -17
rect -190 -119 -156 -85
rect -190 -187 -156 -153
rect -190 -255 -156 -221
rect -190 -323 -156 -289
rect -190 -391 -156 -357
rect -190 -459 -156 -425
rect -190 -527 -156 -493
rect -190 -595 -156 -561
rect 156 561 190 595
rect 156 493 190 527
rect 156 425 190 459
rect 156 357 190 391
rect 156 289 190 323
rect 156 221 190 255
rect 156 153 190 187
rect 156 85 190 119
rect 156 17 190 51
rect 156 -51 190 -17
rect 156 -119 190 -85
rect 156 -187 190 -153
rect 156 -255 190 -221
rect 156 -323 190 -289
rect 156 -391 190 -357
rect 156 -459 190 -425
rect 156 -527 190 -493
rect 156 -595 190 -561
rect -190 -663 -156 -629
rect 156 -663 190 -629
rect -85 -783 -51 -749
rect -17 -783 17 -749
rect 51 -783 85 -749
<< poly >>
rect -33 681 33 697
rect -33 647 -17 681
rect 17 647 33 681
rect -33 631 33 647
rect -30 600 30 631
rect -30 -631 30 -600
rect -33 -647 33 -631
rect -33 -681 -17 -647
rect 17 -681 33 -647
rect -33 -697 33 -681
<< polycont >>
rect -17 647 17 681
rect -17 -681 17 -647
<< locali >>
rect -190 749 -85 783
rect -51 749 -17 783
rect 17 749 51 783
rect 85 749 190 783
rect -190 663 -156 749
rect -33 647 -17 681
rect 17 647 33 681
rect 156 663 190 749
rect -190 595 -156 629
rect -190 527 -156 561
rect -190 459 -156 493
rect -190 391 -156 425
rect -190 323 -156 357
rect -190 255 -156 289
rect -190 187 -156 221
rect -190 119 -156 153
rect -190 51 -156 85
rect -190 -17 -156 17
rect -190 -85 -156 -51
rect -190 -153 -156 -119
rect -190 -221 -156 -187
rect -190 -289 -156 -255
rect -190 -357 -156 -323
rect -190 -425 -156 -391
rect -190 -493 -156 -459
rect -190 -561 -156 -527
rect -190 -629 -156 -595
rect -76 561 -42 604
rect -76 493 -42 523
rect -76 425 -42 451
rect -76 357 -42 379
rect -76 289 -42 307
rect -76 221 -42 235
rect -76 153 -42 163
rect -76 85 -42 91
rect -76 17 -42 19
rect -76 -19 -42 -17
rect -76 -91 -42 -85
rect -76 -163 -42 -153
rect -76 -235 -42 -221
rect -76 -307 -42 -289
rect -76 -379 -42 -357
rect -76 -451 -42 -425
rect -76 -523 -42 -493
rect -76 -604 -42 -561
rect 42 561 76 604
rect 42 493 76 523
rect 42 425 76 451
rect 42 357 76 379
rect 42 289 76 307
rect 42 221 76 235
rect 42 153 76 163
rect 42 85 76 91
rect 42 17 76 19
rect 42 -19 76 -17
rect 42 -91 76 -85
rect 42 -163 76 -153
rect 42 -235 76 -221
rect 42 -307 76 -289
rect 42 -379 76 -357
rect 42 -451 76 -425
rect 42 -523 76 -493
rect 42 -604 76 -561
rect 156 595 190 629
rect 156 527 190 561
rect 156 459 190 493
rect 156 391 190 425
rect 156 323 190 357
rect 156 255 190 289
rect 156 187 190 221
rect 156 119 190 153
rect 156 51 190 85
rect 156 -17 190 17
rect 156 -85 190 -51
rect 156 -153 190 -119
rect 156 -221 190 -187
rect 156 -289 190 -255
rect 156 -357 190 -323
rect 156 -425 190 -391
rect 156 -493 190 -459
rect 156 -561 190 -527
rect 156 -629 190 -595
rect -190 -749 -156 -663
rect -33 -681 -17 -647
rect 17 -681 33 -647
rect 156 -749 190 -663
rect -190 -783 -85 -749
rect -51 -783 -17 -749
rect 17 -783 51 -749
rect 85 -783 190 -749
<< viali >>
rect -17 647 17 681
rect -76 527 -42 557
rect -76 523 -42 527
rect -76 459 -42 485
rect -76 451 -42 459
rect -76 391 -42 413
rect -76 379 -42 391
rect -76 323 -42 341
rect -76 307 -42 323
rect -76 255 -42 269
rect -76 235 -42 255
rect -76 187 -42 197
rect -76 163 -42 187
rect -76 119 -42 125
rect -76 91 -42 119
rect -76 51 -42 53
rect -76 19 -42 51
rect -76 -51 -42 -19
rect -76 -53 -42 -51
rect -76 -119 -42 -91
rect -76 -125 -42 -119
rect -76 -187 -42 -163
rect -76 -197 -42 -187
rect -76 -255 -42 -235
rect -76 -269 -42 -255
rect -76 -323 -42 -307
rect -76 -341 -42 -323
rect -76 -391 -42 -379
rect -76 -413 -42 -391
rect -76 -459 -42 -451
rect -76 -485 -42 -459
rect -76 -527 -42 -523
rect -76 -557 -42 -527
rect 42 527 76 557
rect 42 523 76 527
rect 42 459 76 485
rect 42 451 76 459
rect 42 391 76 413
rect 42 379 76 391
rect 42 323 76 341
rect 42 307 76 323
rect 42 255 76 269
rect 42 235 76 255
rect 42 187 76 197
rect 42 163 76 187
rect 42 119 76 125
rect 42 91 76 119
rect 42 51 76 53
rect 42 19 76 51
rect 42 -51 76 -19
rect 42 -53 76 -51
rect 42 -119 76 -91
rect 42 -125 76 -119
rect 42 -187 76 -163
rect 42 -197 76 -187
rect 42 -255 76 -235
rect 42 -269 76 -255
rect 42 -323 76 -307
rect 42 -341 76 -323
rect 42 -391 76 -379
rect 42 -413 76 -391
rect 42 -459 76 -451
rect 42 -485 76 -459
rect 42 -527 76 -523
rect 42 -557 76 -527
rect -17 -681 17 -647
<< metal1 >>
rect -29 681 29 687
rect -29 647 -17 681
rect 17 647 29 681
rect -29 641 29 647
rect -82 557 -36 600
rect -82 523 -76 557
rect -42 523 -36 557
rect -82 485 -36 523
rect -82 451 -76 485
rect -42 451 -36 485
rect -82 413 -36 451
rect -82 379 -76 413
rect -42 379 -36 413
rect -82 341 -36 379
rect -82 307 -76 341
rect -42 307 -36 341
rect -82 269 -36 307
rect -82 235 -76 269
rect -42 235 -36 269
rect -82 197 -36 235
rect -82 163 -76 197
rect -42 163 -36 197
rect -82 125 -36 163
rect -82 91 -76 125
rect -42 91 -36 125
rect -82 53 -36 91
rect -82 19 -76 53
rect -42 19 -36 53
rect -82 -19 -36 19
rect -82 -53 -76 -19
rect -42 -53 -36 -19
rect -82 -91 -36 -53
rect -82 -125 -76 -91
rect -42 -125 -36 -91
rect -82 -163 -36 -125
rect -82 -197 -76 -163
rect -42 -197 -36 -163
rect -82 -235 -36 -197
rect -82 -269 -76 -235
rect -42 -269 -36 -235
rect -82 -307 -36 -269
rect -82 -341 -76 -307
rect -42 -341 -36 -307
rect -82 -379 -36 -341
rect -82 -413 -76 -379
rect -42 -413 -36 -379
rect -82 -451 -36 -413
rect -82 -485 -76 -451
rect -42 -485 -36 -451
rect -82 -523 -36 -485
rect -82 -557 -76 -523
rect -42 -557 -36 -523
rect -82 -600 -36 -557
rect 36 557 82 600
rect 36 523 42 557
rect 76 523 82 557
rect 36 485 82 523
rect 36 451 42 485
rect 76 451 82 485
rect 36 413 82 451
rect 36 379 42 413
rect 76 379 82 413
rect 36 341 82 379
rect 36 307 42 341
rect 76 307 82 341
rect 36 269 82 307
rect 36 235 42 269
rect 76 235 82 269
rect 36 197 82 235
rect 36 163 42 197
rect 76 163 82 197
rect 36 125 82 163
rect 36 91 42 125
rect 76 91 82 125
rect 36 53 82 91
rect 36 19 42 53
rect 76 19 82 53
rect 36 -19 82 19
rect 36 -53 42 -19
rect 76 -53 82 -19
rect 36 -91 82 -53
rect 36 -125 42 -91
rect 76 -125 82 -91
rect 36 -163 82 -125
rect 36 -197 42 -163
rect 76 -197 82 -163
rect 36 -235 82 -197
rect 36 -269 42 -235
rect 76 -269 82 -235
rect 36 -307 82 -269
rect 36 -341 42 -307
rect 76 -341 82 -307
rect 36 -379 82 -341
rect 36 -413 42 -379
rect 76 -413 82 -379
rect 36 -451 82 -413
rect 36 -485 42 -451
rect 76 -485 82 -451
rect 36 -523 82 -485
rect 36 -557 42 -523
rect 76 -557 82 -523
rect 36 -600 82 -557
rect -29 -647 29 -641
rect -29 -681 -17 -647
rect 17 -681 29 -647
rect -29 -687 29 -681
<< properties >>
string FIXED_BBOX -173 -766 173 766
<< end >>
