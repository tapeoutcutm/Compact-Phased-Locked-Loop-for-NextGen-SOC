magic
tech sky130A
magscale 1 2
timestamp 1713524523
<< nwell >>
rect 6072 16 6320 306
rect 4908 -654 5156 -364
rect 5498 -1322 5746 -1032
<< pwell >>
rect 6062 -262 6198 -64
rect 4838 -948 4974 -750
rect 5496 -1598 5632 -1400
<< psubdiff >>
rect 6088 -141 6172 -90
rect 6088 -175 6114 -141
rect 6148 -175 6172 -141
rect 6088 -236 6172 -175
rect 4864 -827 4948 -776
rect 4864 -861 4890 -827
rect 4924 -861 4948 -827
rect 4864 -922 4948 -861
rect 5522 -1477 5606 -1426
rect 5522 -1511 5548 -1477
rect 5582 -1511 5606 -1477
rect 5522 -1572 5606 -1511
<< nsubdiff >>
rect 6108 210 6274 260
rect 6108 176 6174 210
rect 6208 176 6274 210
rect 6108 142 6274 176
rect 6108 108 6174 142
rect 6208 108 6274 142
rect 6108 66 6274 108
rect 4944 -460 5110 -410
rect 4944 -494 5010 -460
rect 5044 -494 5110 -460
rect 4944 -528 5110 -494
rect 4944 -562 5010 -528
rect 5044 -562 5110 -528
rect 4944 -604 5110 -562
rect 5534 -1128 5700 -1078
rect 5534 -1162 5600 -1128
rect 5634 -1162 5700 -1128
rect 5534 -1196 5700 -1162
rect 5534 -1230 5600 -1196
rect 5634 -1230 5700 -1196
rect 5534 -1272 5700 -1230
<< psubdiffcont >>
rect 6114 -175 6148 -141
rect 4890 -861 4924 -827
rect 5548 -1511 5582 -1477
<< nsubdiffcont >>
rect 6174 176 6208 210
rect 6174 108 6208 142
rect 5010 -494 5044 -460
rect 5010 -562 5044 -528
rect 5600 -1162 5634 -1128
rect 5600 -1230 5634 -1196
<< locali >>
rect 2500 204 2538 262
rect 6034 248 6274 290
rect 6108 210 6274 248
rect 6108 176 6174 210
rect 6208 176 6274 210
rect 6108 142 6274 176
rect 6108 108 6174 142
rect 6208 108 6274 142
rect 6108 66 6274 108
rect 6006 -11 6056 20
rect 2158 -31 2280 -20
rect 2158 -65 2166 -31
rect 2200 -65 2238 -31
rect 2272 -65 2280 -31
rect 2158 -76 2280 -65
rect 4060 -26 4108 -14
rect 4060 -60 4067 -26
rect 4101 -60 4108 -26
rect 4536 -23 4570 -22
rect 4536 -58 4570 -57
rect 4896 -60 5068 -14
rect 5436 -60 5608 -14
rect 6006 -45 6014 -11
rect 6048 -45 6056 -11
rect 4060 -72 4108 -60
rect 6006 -76 6056 -45
rect 6088 -141 6172 -90
rect 6088 -175 6114 -141
rect 6148 -175 6172 -141
rect 6088 -256 6172 -175
rect 6004 -272 6172 -256
rect 6034 -294 6172 -272
rect 4870 -420 5110 -380
rect 4944 -460 5110 -420
rect 4944 -494 5010 -460
rect 5044 -494 5110 -460
rect 4944 -528 5110 -494
rect 4944 -562 5010 -528
rect 5044 -562 5110 -528
rect 4944 -604 5110 -562
rect 3808 -674 3858 -644
rect 3808 -708 3816 -674
rect 3850 -708 3858 -674
rect 3808 -738 3858 -708
rect 4220 -732 4428 -682
rect 4614 -718 4622 -684
rect 4656 -718 4664 -684
rect 4752 -716 4760 -682
rect 4794 -716 4802 -682
rect 4864 -827 4948 -776
rect 4864 -861 4890 -827
rect 4924 -861 4948 -827
rect 4864 -928 4948 -861
rect 4620 -930 4948 -928
rect 4864 -962 4948 -930
rect 2502 -1124 2540 -1084
rect 5460 -1088 5700 -1050
rect 5534 -1128 5700 -1088
rect 5534 -1162 5600 -1128
rect 5634 -1162 5700 -1128
rect 5534 -1196 5700 -1162
rect 5534 -1230 5600 -1196
rect 5634 -1230 5700 -1196
rect 5534 -1272 5700 -1230
rect 5428 -1343 5492 -1310
rect 2236 -1360 2284 -1350
rect 4496 -1355 4530 -1354
rect 2236 -1394 2243 -1360
rect 2277 -1394 2284 -1360
rect 2236 -1404 2284 -1394
rect 4068 -1362 4102 -1356
rect 4496 -1390 4530 -1389
rect 4068 -1402 4102 -1396
rect 4846 -1398 5024 -1350
rect 5428 -1377 5443 -1343
rect 5477 -1377 5492 -1343
rect 5428 -1410 5492 -1377
rect 5522 -1477 5606 -1426
rect 5522 -1511 5548 -1477
rect 5582 -1511 5606 -1477
rect 5522 -1594 5606 -1511
rect 5428 -1600 5606 -1594
rect 5458 -1630 5606 -1600
<< viali >>
rect 2166 -65 2200 -31
rect 2238 -65 2272 -31
rect 4067 -60 4101 -26
rect 4536 -57 4570 -23
rect 6014 -45 6048 -11
rect 3816 -708 3850 -674
rect 4622 -718 4656 -684
rect 4760 -716 4794 -682
rect 2243 -1394 2277 -1360
rect 4068 -1396 4102 -1362
rect 4496 -1389 4530 -1355
rect 5443 -1377 5477 -1343
<< metal1 >>
rect 1912 314 2112 514
rect 1912 218 2224 314
rect 4132 220 4540 314
rect 4962 218 5318 314
rect 5498 218 5574 314
rect 5750 218 6104 314
rect 1572 38 1772 78
rect 1572 -14 1680 38
rect 1732 -14 1772 38
rect 1572 -26 1772 -14
rect 1572 -78 1680 -26
rect 1732 -78 1772 -26
rect 1572 -122 1772 -78
rect 1912 -354 2044 218
rect 6366 32 6566 88
rect 3644 -2 3730 0
rect 2146 -22 2292 -14
rect 2146 -74 2161 -22
rect 2213 -74 2225 -22
rect 2277 -74 2292 -22
rect 3644 -54 3661 -2
rect 3713 -54 3730 -2
rect 4054 -12 4114 -2
rect 3644 -56 3730 -54
rect 4040 -17 4128 -12
rect 4040 -69 4058 -17
rect 4110 -69 4128 -17
rect 4040 -74 4128 -69
rect 4514 -13 4586 -6
rect 4514 -65 4524 -13
rect 4576 -65 4586 -13
rect 4514 -72 4586 -65
rect 6000 -11 6566 32
rect 6000 -45 6014 -11
rect 6048 -45 6566 -11
rect 2146 -82 2292 -74
rect 4054 -84 4114 -74
rect 6000 -88 6566 -45
rect 6366 -112 6566 -88
rect 4132 -326 4504 -230
rect 4962 -326 5574 -230
rect 5652 -326 6306 -230
rect 1912 -450 3782 -354
rect 4242 -450 4318 -354
rect 1912 -1022 2044 -450
rect 3802 -640 3864 -632
rect 3728 -664 3864 -640
rect 3728 -716 3738 -664
rect 3790 -716 3802 -664
rect 3854 -716 3864 -664
rect 4592 -673 4680 -668
rect 3728 -740 3864 -716
rect 4220 -732 4434 -680
rect 4592 -725 4610 -673
rect 4662 -725 4680 -673
rect 4592 -730 4680 -725
rect 4732 -673 4820 -668
rect 4732 -725 4750 -673
rect 4802 -725 4820 -673
rect 4732 -730 4820 -725
rect 3802 -750 3864 -740
rect 6174 -898 6306 -326
rect 3782 -994 6306 -898
rect 1912 -1118 2226 -1022
rect 4132 -1116 5652 -1022
rect 1572 -1318 1772 -1288
rect 5422 -1302 5698 -1298
rect 1572 -1334 1782 -1318
rect 1572 -1386 1704 -1334
rect 1756 -1386 1782 -1334
rect 3644 -1334 3730 -1332
rect 1572 -1398 1782 -1386
rect 1572 -1450 1704 -1398
rect 1756 -1450 1782 -1398
rect 2210 -1350 2300 -1336
rect 2210 -1402 2229 -1350
rect 2281 -1402 2300 -1350
rect 3644 -1386 3661 -1334
rect 3713 -1386 3730 -1334
rect 4062 -1348 4108 -1344
rect 3644 -1388 3730 -1386
rect 4040 -1353 4128 -1348
rect 4490 -1352 4536 -1342
rect 5422 -1343 5509 -1302
rect 2210 -1416 2300 -1402
rect 4040 -1405 4058 -1353
rect 4110 -1405 4128 -1353
rect 4040 -1410 4128 -1405
rect 4476 -1355 4548 -1352
rect 4476 -1357 4496 -1355
rect 4530 -1357 4548 -1355
rect 4476 -1409 4486 -1357
rect 4538 -1409 4548 -1357
rect 4062 -1414 4108 -1410
rect 4476 -1414 4548 -1409
rect 5422 -1377 5443 -1343
rect 5477 -1354 5509 -1343
rect 5561 -1354 5698 -1302
rect 5477 -1366 5698 -1354
rect 5477 -1377 5509 -1366
rect 5422 -1418 5509 -1377
rect 5561 -1418 5698 -1366
rect 5422 -1422 5584 -1418
rect 1572 -1466 1782 -1450
rect 1572 -1488 1772 -1466
rect 6174 -1566 6306 -994
rect 6366 -1298 6566 -1262
rect 6356 -1300 6566 -1298
rect 6356 -1352 6375 -1300
rect 6427 -1352 6566 -1300
rect 6356 -1364 6566 -1352
rect 6356 -1416 6375 -1364
rect 6427 -1416 6566 -1364
rect 6356 -1418 6566 -1416
rect 6366 -1462 6566 -1418
rect 4132 -1662 6306 -1566
rect 6106 -1860 6306 -1662
<< via1 >>
rect 1680 -14 1732 38
rect 1680 -78 1732 -26
rect 2161 -31 2213 -22
rect 2161 -65 2166 -31
rect 2166 -65 2200 -31
rect 2200 -65 2213 -31
rect 2161 -74 2213 -65
rect 2225 -31 2277 -22
rect 2225 -65 2238 -31
rect 2238 -65 2272 -31
rect 2272 -65 2277 -31
rect 2225 -74 2277 -65
rect 3661 -54 3713 -2
rect 4058 -26 4110 -17
rect 4058 -60 4067 -26
rect 4067 -60 4101 -26
rect 4101 -60 4110 -26
rect 4058 -69 4110 -60
rect 4524 -23 4576 -13
rect 4524 -57 4536 -23
rect 4536 -57 4570 -23
rect 4570 -57 4576 -23
rect 4524 -65 4576 -57
rect 3738 -716 3790 -664
rect 3802 -674 3854 -664
rect 3802 -708 3816 -674
rect 3816 -708 3850 -674
rect 3850 -708 3854 -674
rect 3802 -716 3854 -708
rect 4610 -684 4662 -673
rect 4610 -718 4622 -684
rect 4622 -718 4656 -684
rect 4656 -718 4662 -684
rect 4610 -725 4662 -718
rect 4750 -682 4802 -673
rect 4750 -716 4760 -682
rect 4760 -716 4794 -682
rect 4794 -716 4802 -682
rect 4750 -725 4802 -716
rect 1704 -1386 1756 -1334
rect 1704 -1450 1756 -1398
rect 2229 -1360 2281 -1350
rect 2229 -1394 2243 -1360
rect 2243 -1394 2277 -1360
rect 2277 -1394 2281 -1360
rect 2229 -1402 2281 -1394
rect 3661 -1386 3713 -1334
rect 4058 -1362 4110 -1353
rect 4058 -1396 4068 -1362
rect 4068 -1396 4102 -1362
rect 4102 -1396 4110 -1362
rect 4058 -1405 4110 -1396
rect 4486 -1389 4496 -1357
rect 4496 -1389 4530 -1357
rect 4530 -1389 4538 -1357
rect 4486 -1409 4538 -1389
rect 5509 -1354 5561 -1302
rect 5509 -1418 5561 -1366
rect 6375 -1352 6427 -1300
rect 6375 -1416 6427 -1364
<< metal2 >>
rect 1744 54 2281 60
rect 1664 38 2281 54
rect 1664 -14 1680 38
rect 1732 -14 2281 38
rect 1664 -22 2281 -14
rect 1664 -26 2161 -22
rect 1664 -78 1680 -26
rect 1732 -74 2161 -26
rect 2213 -74 2225 -22
rect 2277 -74 2281 -22
rect 1732 -78 2281 -74
rect 1664 -94 2281 -78
rect 3654 -2 3720 10
rect 3654 -54 3661 -2
rect 3713 -54 3720 -2
rect 3654 -630 3720 -54
rect 4050 -13 4584 6
rect 4050 -17 4524 -13
rect 4050 -69 4058 -17
rect 4110 -65 4524 -17
rect 4576 -65 4584 -13
rect 4110 -69 4584 -65
rect 4050 -82 4584 -69
rect 4050 -506 4118 -82
rect 4050 -564 4810 -506
rect 3654 -664 3854 -630
rect 3654 -716 3738 -664
rect 3790 -716 3802 -664
rect 4602 -673 4670 -658
rect 4602 -674 4610 -673
rect 3654 -750 3854 -716
rect 4050 -725 4610 -674
rect 4662 -725 4670 -673
rect 4050 -732 4670 -725
rect 1674 -1334 2308 -1310
rect 1674 -1386 1704 -1334
rect 1756 -1350 2308 -1334
rect 1756 -1386 2229 -1350
rect 1674 -1398 2229 -1386
rect 1674 -1450 1704 -1398
rect 1756 -1402 2229 -1398
rect 2281 -1402 2308 -1350
rect 3654 -1334 3720 -750
rect 3654 -1386 3661 -1334
rect 3713 -1386 3720 -1334
rect 3654 -1398 3720 -1386
rect 4050 -1340 4118 -732
rect 4602 -740 4670 -732
rect 4742 -673 4810 -564
rect 4742 -725 4750 -673
rect 4802 -725 4810 -673
rect 4742 -740 4810 -725
rect 5496 -1298 5574 -1288
rect 6366 -1298 6436 -1288
rect 5496 -1300 6436 -1298
rect 5496 -1302 6375 -1300
rect 4050 -1353 4544 -1340
rect 1756 -1450 2308 -1402
rect 4050 -1405 4058 -1353
rect 4110 -1357 4544 -1353
rect 4110 -1405 4486 -1357
rect 4050 -1409 4486 -1405
rect 4538 -1409 4544 -1357
rect 4050 -1424 4544 -1409
rect 5496 -1354 5509 -1302
rect 5561 -1352 6375 -1302
rect 6427 -1352 6436 -1300
rect 5561 -1354 6436 -1352
rect 5496 -1364 6436 -1354
rect 5496 -1366 6375 -1364
rect 5496 -1418 5509 -1366
rect 5561 -1416 6375 -1366
rect 6427 -1416 6436 -1364
rect 5561 -1418 6436 -1416
rect 5496 -1432 5574 -1418
rect 6366 -1428 6436 -1418
rect 1674 -1460 2308 -1450
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1712078602
transform 1 0 2126 0 1 -1614
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_1
timestamp 1712078602
transform 1 0 2126 0 1 -278
box -38 -48 130 592
use sky130_fd_sc_hd__dfrbp_2#0  x1
timestamp 1712816020
transform 1 0 2218 0 1 -278
box -38 -48 2246 592
use sky130_fd_sc_hd__dfrbp_2#0  x2
timestamp 1712816020
transform 1 0 2218 0 1 -1614
box -38 -48 2246 592
use sky130_fd_sc_hd__and2_2#0  x3
timestamp 1712816020
transform -1 0 4870 0 1 -946
box -38 -48 590 592
use sky130_fd_sc_hd__inv_4#0  x4
timestamp 1712816020
transform -1 0 4242 0 1 -946
box -38 -48 498 592
use sky130_fd_sc_hd__inv_4#0  x5
timestamp 1712816020
transform 1 0 4464 0 1 -1614
box -38 -48 498 592
use sky130_fd_sc_hd__inv_4#0  x6
timestamp 1712816020
transform 1 0 5000 0 1 -1614
box -38 -48 498 592
use sky130_fd_sc_hd__inv_4#0  x7
timestamp 1712816020
transform 1 0 4502 0 1 -278
box -38 -48 498 592
use sky130_fd_sc_hd__inv_4#0  x8
timestamp 1712816020
transform 1 0 5038 0 1 -278
box -38 -48 498 592
use sky130_fd_sc_hd__inv_4#0  x9
timestamp 1712816020
transform 1 0 5574 0 1 -278
box -38 -48 498 592
<< labels >>
flabel metal1 s 6366 -112 6566 88 0 FreeSans 626 0 0 0 QA
port 1 nsew
flabel metal1 s 1572 -122 1772 78 0 FreeSans 626 0 0 0 A
port 2 nsew
flabel metal1 s 1912 314 2112 514 0 FreeSans 626 180 0 0 VDD
port 3 nsew
flabel metal1 s 6106 -1860 6306 -1660 0 FreeSans 626 180 0 0 VSS
port 4 nsew
flabel metal1 s 1572 -1488 1772 -1288 0 FreeSans 626 0 0 0 B
port 5 nsew
flabel metal1 s 6366 -1462 6566 -1262 0 FreeSans 626 0 0 0 QB
port 6 nsew
<< end >>
