VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_vks_pll
  CLASS BLOCK ;
  FOREIGN tt_um_vks_pll ;
  ORIGIN 0.000 0.000 ;
  SIZE 334.880 BY 225.760 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 154.870 224.760 155.170 225.760 ;
    END
  END clk
  PIN ena
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 158.550 224.760 158.850 225.760 ;
    END
  END ena
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 151.190 224.760 151.490 225.760 ;
    END
  END rst_n
  PIN ua[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met4 ;
        RECT 156.560 0.000 157.160 1.000 ;
    END
  END ua[0]
  PIN ua[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met4 ;
        RECT 134.480 0.000 135.080 1.000 ;
    END
  END ua[1]
  PIN ua[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.511500 ;
    PORT
      LAYER met4 ;
        RECT 112.400 0.000 113.000 1.000 ;
    END
  END ua[2]
  PIN ua[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.511500 ;
    PORT
      LAYER met4 ;
        RECT 90.320 0.000 90.920 1.000 ;
    END
  END ua[3]
  PIN ua[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 68.240 0.000 68.840 1.000 ;
    END
  END ua[4]
  PIN ua[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 46.160 0.000 46.760 1.000 ;
    END
  END ua[5]
  PIN ua[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 24.080 0.000 24.680 1.000 ;
    END
  END ua[6]
  PIN ua[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 2.000 0.000 2.600 1.000 ;
    END
  END ua[7]
  PIN ui_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 147.510 224.760 147.810 225.760 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 143.830 224.760 144.130 225.760 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 140.150 224.760 140.450 225.760 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 136.470 224.760 136.770 225.760 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 132.790 224.760 133.090 225.760 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 129.110 224.760 129.410 225.760 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 125.430 224.760 125.730 225.760 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 121.750 224.760 122.050 225.760 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 118.070 224.760 118.370 225.760 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 114.390 224.760 114.690 225.760 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 110.710 224.760 111.010 225.760 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 107.030 224.760 107.330 225.760 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 103.350 224.760 103.650 225.760 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 99.670 224.760 99.970 225.760 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 95.990 224.760 96.290 225.760 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 92.310 224.760 92.610 225.760 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 29.750 224.760 30.050 225.760 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 26.070 224.760 26.370 225.760 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 22.390 224.760 22.690 225.760 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 18.710 224.760 19.010 225.760 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 15.030 224.760 15.330 225.760 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 11.350 224.760 11.650 225.760 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 7.670 224.760 7.970 225.760 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 3.990 224.760 4.290 225.760 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 59.190 224.760 59.490 225.760 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 55.510 224.760 55.810 225.760 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 51.830 224.760 52.130 225.760 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 48.150 224.760 48.450 225.760 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 44.470 224.760 44.770 225.760 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 40.790 224.760 41.090 225.760 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 37.110 224.760 37.410 225.760 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 33.430 224.760 33.730 225.760 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 88.630 224.760 88.930 225.760 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 84.950 224.760 85.250 225.760 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 81.270 224.760 81.570 225.760 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 77.590 224.760 77.890 225.760 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 73.910 224.760 74.210 225.760 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 70.230 224.760 70.530 225.760 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 66.550 224.760 66.850 225.760 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 62.870 224.760 63.170 225.760 ;
    END
  END uo_out[7]
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1.000 5.000 2.500 220.760 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 49.000 5.000 50.500 220.760 ;
    END
  END VGND
  OBS
      LAYER nwell ;
        RECT 115.420 23.230 116.440 23.280 ;
        RECT 115.420 23.190 116.600 23.230 ;
        RECT 115.420 21.585 127.760 23.190 ;
        RECT 115.420 21.580 116.440 21.585 ;
      LAYER pwell ;
        RECT 116.640 21.290 118.920 21.295 ;
        RECT 115.490 21.065 118.920 21.290 ;
        RECT 122.125 21.065 123.055 21.285 ;
        RECT 115.490 20.610 127.565 21.065 ;
        RECT 116.640 20.385 127.565 20.610 ;
        RECT 127.255 20.195 127.425 20.385 ;
      LAYER nwell ;
        RECT 116.800 19.490 117.830 19.510 ;
        RECT 120.800 19.490 123.080 19.500 ;
        RECT 116.800 19.440 123.080 19.490 ;
        RECT 116.800 17.885 125.590 19.440 ;
        RECT 116.800 17.880 117.830 17.885 ;
        RECT 120.800 17.850 125.590 17.885 ;
        RECT 122.910 17.835 125.590 17.850 ;
      LAYER pwell ;
        RECT 116.910 17.505 118.120 17.560 ;
        RECT 119.085 17.550 120.675 17.595 ;
        RECT 119.085 17.545 123.160 17.550 ;
        RECT 119.085 17.505 125.345 17.545 ;
        RECT 116.910 16.900 125.345 17.505 ;
        RECT 118.105 16.690 125.345 16.900 ;
        RECT 118.105 16.685 120.675 16.690 ;
        RECT 118.105 16.665 118.245 16.685 ;
        RECT 118.075 16.495 118.245 16.665 ;
        RECT 123.155 16.635 125.345 16.690 ;
        RECT 123.245 16.445 123.415 16.635 ;
      LAYER nwell ;
        RECT 115.670 14.190 127.990 15.780 ;
        RECT 116.570 14.175 127.990 14.190 ;
      LAYER pwell ;
        RECT 115.790 13.885 116.910 13.960 ;
        RECT 115.790 13.655 119.150 13.885 ;
        RECT 122.355 13.655 123.285 13.875 ;
        RECT 115.790 12.990 127.795 13.655 ;
        RECT 116.870 12.975 127.795 12.990 ;
        RECT 127.485 12.785 127.655 12.975 ;
      LAYER li1 ;
        RECT 116.100 23.085 116.670 23.090 ;
        RECT 116.100 22.920 127.570 23.085 ;
        RECT 116.105 22.340 116.275 22.920 ;
        RECT 116.530 22.915 127.570 22.920 ;
        RECT 116.810 21.725 116.980 22.915 ;
        RECT 117.150 22.360 117.450 22.745 ;
        RECT 117.620 22.535 117.950 22.915 ;
        RECT 118.500 22.485 118.840 22.915 ;
        RECT 117.150 21.815 117.540 22.360 ;
        RECT 119.010 22.315 119.235 22.745 ;
        RECT 119.515 22.535 119.860 22.915 ;
        RECT 120.040 22.365 120.210 22.655 ;
        RECT 120.380 22.455 120.630 22.915 ;
        RECT 117.735 22.145 119.235 22.315 ;
        RECT 115.530 21.120 116.450 21.270 ;
        RECT 115.530 20.630 116.470 21.120 ;
        RECT 115.530 20.620 116.450 20.630 ;
        RECT 116.810 20.365 116.980 21.210 ;
        RECT 117.150 21.105 117.320 21.815 ;
        RECT 117.735 21.605 117.905 22.145 ;
        RECT 118.580 22.075 119.235 22.145 ;
        RECT 119.410 22.195 120.210 22.365 ;
        RECT 120.800 22.405 121.670 22.745 ;
        RECT 117.490 21.275 117.905 21.605 ;
        RECT 117.150 20.590 117.530 21.105 ;
        RECT 117.700 20.365 117.870 21.105 ;
        RECT 118.075 20.545 118.410 21.975 ;
        RECT 118.580 21.165 118.750 22.075 ;
        RECT 119.410 21.605 119.580 22.195 ;
        RECT 120.800 22.025 120.970 22.405 ;
        RECT 121.905 22.285 122.075 22.745 ;
        RECT 122.245 22.455 122.615 22.915 ;
        RECT 122.910 22.315 123.080 22.655 ;
        RECT 123.250 22.485 123.580 22.915 ;
        RECT 123.815 22.315 123.985 22.655 ;
        RECT 119.750 21.855 120.970 22.025 ;
        RECT 121.140 21.945 121.600 22.235 ;
        RECT 121.905 22.115 122.465 22.285 ;
        RECT 122.910 22.145 123.985 22.315 ;
        RECT 124.155 22.415 124.835 22.745 ;
        RECT 125.050 22.415 125.300 22.745 ;
        RECT 125.470 22.455 125.720 22.915 ;
        RECT 125.890 22.730 126.210 22.915 ;
        RECT 122.295 21.975 122.465 22.115 ;
        RECT 121.140 21.935 122.105 21.945 ;
        RECT 120.800 21.765 120.970 21.855 ;
        RECT 121.430 21.775 122.105 21.935 ;
        RECT 118.920 21.575 119.580 21.605 ;
        RECT 118.920 21.355 119.755 21.575 ;
        RECT 119.410 21.275 119.755 21.355 ;
        RECT 118.580 20.995 119.235 21.165 ;
        RECT 118.580 20.365 118.815 20.825 ;
        RECT 118.985 20.625 119.235 20.995 ;
        RECT 119.585 20.745 119.755 21.275 ;
        RECT 119.925 21.315 120.465 21.685 ;
        RECT 120.800 21.595 121.205 21.765 ;
        RECT 119.925 20.915 120.165 21.315 ;
        RECT 120.645 21.145 120.865 21.425 ;
        RECT 120.335 20.975 120.865 21.145 ;
        RECT 120.335 20.745 120.505 20.975 ;
        RECT 121.035 20.815 121.205 21.595 ;
        RECT 121.375 20.985 121.725 21.605 ;
        RECT 121.895 20.985 122.105 21.775 ;
        RECT 122.295 21.805 123.795 21.975 ;
        RECT 122.295 21.115 122.465 21.805 ;
        RECT 124.155 21.635 124.325 22.415 ;
        RECT 125.130 22.285 125.300 22.415 ;
        RECT 122.635 21.465 124.325 21.635 ;
        RECT 124.495 21.855 124.960 22.245 ;
        RECT 125.130 22.115 125.525 22.285 ;
        RECT 122.635 21.285 122.805 21.465 ;
        RECT 119.585 20.575 120.505 20.745 ;
        RECT 120.675 20.365 120.865 20.805 ;
        RECT 121.035 20.535 121.985 20.815 ;
        RECT 122.295 20.725 122.555 21.115 ;
        RECT 122.975 21.045 123.765 21.295 ;
        RECT 122.205 20.555 122.555 20.725 ;
        RECT 122.765 20.365 123.095 20.825 ;
        RECT 123.970 20.755 124.140 21.465 ;
        RECT 124.495 21.265 124.665 21.855 ;
        RECT 124.310 21.045 124.665 21.265 ;
        RECT 124.835 21.045 125.185 21.665 ;
        RECT 125.355 20.755 125.525 22.115 ;
        RECT 125.890 21.945 126.215 22.730 ;
        RECT 125.695 20.895 126.155 21.945 ;
        RECT 123.970 20.585 124.825 20.755 ;
        RECT 125.030 20.585 125.525 20.755 ;
        RECT 125.695 20.365 126.025 20.725 ;
        RECT 126.385 20.625 126.555 22.745 ;
        RECT 126.725 22.415 127.055 22.915 ;
        RECT 127.225 22.245 127.480 22.745 ;
        RECT 126.730 22.075 127.480 22.245 ;
        RECT 126.730 21.085 126.960 22.075 ;
        RECT 127.130 21.890 127.480 21.905 ;
        RECT 127.130 21.880 130.510 21.890 ;
        RECT 127.130 21.280 131.200 21.880 ;
        RECT 127.130 21.255 127.480 21.280 ;
        RECT 130.250 21.270 131.200 21.280 ;
        RECT 126.730 20.915 127.480 21.085 ;
        RECT 126.725 20.365 127.055 20.745 ;
        RECT 127.225 20.625 127.480 20.915 ;
        RECT 116.530 20.195 127.570 20.365 ;
        RECT 117.170 19.385 118.490 19.420 ;
        RECT 117.170 19.215 120.690 19.385 ;
        RECT 117.170 19.210 118.495 19.215 ;
        RECT 117.170 19.180 117.540 19.210 ;
        RECT 117.150 19.010 117.540 19.180 ;
        RECT 113.520 18.230 114.570 18.500 ;
        RECT 117.155 18.430 117.325 19.010 ;
        RECT 118.215 18.545 118.495 19.210 ;
        RECT 118.015 18.230 118.330 18.345 ;
        RECT 113.520 17.905 118.330 18.230 ;
        RECT 118.665 18.325 118.965 18.875 ;
        RECT 119.175 18.495 119.505 19.215 ;
        RECT 119.695 18.495 120.145 19.045 ;
        RECT 118.665 18.155 119.605 18.325 ;
        RECT 118.910 17.905 119.250 17.970 ;
        RECT 119.435 17.905 119.605 18.155 ;
        RECT 113.520 17.670 118.705 17.905 ;
        RECT 113.520 17.610 114.570 17.670 ;
        RECT 118.015 17.655 118.705 17.670 ;
        RECT 118.910 17.660 119.265 17.905 ;
        RECT 118.935 17.655 119.265 17.660 ;
        RECT 119.435 17.575 119.725 17.905 ;
        RECT 119.895 17.900 120.145 18.495 ;
        RECT 120.315 18.075 120.605 19.215 ;
        RECT 123.100 19.165 125.400 19.335 ;
        RECT 123.230 18.025 123.495 19.165 ;
        RECT 123.665 18.195 123.995 18.995 ;
        RECT 124.165 18.365 124.335 19.165 ;
        RECT 124.505 18.215 124.835 18.995 ;
        RECT 125.005 18.705 125.215 19.165 ;
        RECT 124.505 18.195 125.270 18.215 ;
        RECT 123.665 18.050 125.270 18.195 ;
        RECT 125.700 18.050 126.430 18.080 ;
        RECT 123.665 18.025 126.430 18.050 ;
        RECT 120.880 17.900 121.720 17.910 ;
        RECT 119.895 17.850 121.720 17.900 ;
        RECT 123.205 17.850 124.835 17.855 ;
        RECT 119.895 17.640 124.835 17.850 ;
        RECT 119.435 17.485 119.605 17.575 ;
        RECT 116.930 16.930 117.770 17.480 ;
        RECT 118.215 17.295 119.605 17.485 ;
        RECT 118.215 16.935 118.545 17.295 ;
        RECT 119.895 17.125 120.145 17.640 ;
        RECT 120.780 17.630 124.835 17.640 ;
        RECT 120.880 17.605 124.835 17.630 ;
        RECT 120.880 17.600 123.550 17.605 ;
        RECT 120.880 17.590 121.720 17.600 ;
        RECT 119.175 16.665 119.425 17.125 ;
        RECT 119.595 16.835 120.145 17.125 ;
        RECT 120.315 16.665 120.605 17.465 ;
        RECT 125.005 17.460 126.430 18.025 ;
        RECT 125.005 17.435 125.270 17.460 ;
        RECT 123.665 17.255 125.270 17.435 ;
        RECT 125.700 17.410 126.430 17.460 ;
        RECT 117.930 16.495 120.690 16.665 ;
        RECT 123.230 16.615 123.495 17.075 ;
        RECT 123.665 16.785 123.995 17.255 ;
        RECT 124.165 16.615 124.335 17.075 ;
        RECT 124.505 16.785 124.835 17.255 ;
        RECT 125.005 16.615 125.255 17.080 ;
        RECT 123.100 16.445 125.400 16.615 ;
        RECT 116.180 15.675 117.220 15.690 ;
        RECT 116.180 15.505 127.800 15.675 ;
        RECT 116.180 15.500 117.220 15.505 ;
        RECT 116.190 15.470 116.590 15.500 ;
        RECT 116.195 14.890 116.365 15.470 ;
        RECT 117.040 14.315 117.210 15.500 ;
        RECT 117.380 14.950 117.680 15.335 ;
        RECT 117.850 15.125 118.180 15.505 ;
        RECT 118.730 15.075 119.070 15.505 ;
        RECT 117.380 14.405 117.770 14.950 ;
        RECT 119.240 14.905 119.465 15.335 ;
        RECT 119.745 15.125 120.090 15.505 ;
        RECT 120.270 14.955 120.440 15.245 ;
        RECT 120.610 15.045 120.860 15.505 ;
        RECT 117.965 14.735 119.465 14.905 ;
        RECT 115.790 13.750 116.440 13.930 ;
        RECT 115.780 12.840 116.460 13.750 ;
        RECT 117.040 12.955 117.210 13.800 ;
        RECT 117.380 13.695 117.550 14.405 ;
        RECT 117.965 14.195 118.135 14.735 ;
        RECT 118.810 14.665 119.465 14.735 ;
        RECT 119.640 14.785 120.440 14.955 ;
        RECT 121.030 14.995 121.900 15.335 ;
        RECT 117.720 13.865 118.135 14.195 ;
        RECT 117.380 13.180 117.760 13.695 ;
        RECT 117.930 12.955 118.100 13.695 ;
        RECT 118.305 13.135 118.640 14.565 ;
        RECT 118.810 13.755 118.980 14.665 ;
        RECT 119.640 14.195 119.810 14.785 ;
        RECT 121.030 14.615 121.200 14.995 ;
        RECT 122.135 14.875 122.305 15.335 ;
        RECT 122.475 15.045 122.845 15.505 ;
        RECT 123.140 14.905 123.310 15.245 ;
        RECT 123.480 15.075 123.810 15.505 ;
        RECT 124.045 14.905 124.215 15.245 ;
        RECT 119.980 14.445 121.200 14.615 ;
        RECT 121.370 14.535 121.830 14.825 ;
        RECT 122.135 14.705 122.695 14.875 ;
        RECT 123.140 14.735 124.215 14.905 ;
        RECT 124.385 15.005 125.065 15.335 ;
        RECT 125.280 15.005 125.530 15.335 ;
        RECT 125.700 15.045 125.950 15.505 ;
        RECT 126.130 15.320 126.440 15.505 ;
        RECT 122.525 14.565 122.695 14.705 ;
        RECT 121.370 14.525 122.335 14.535 ;
        RECT 121.030 14.355 121.200 14.445 ;
        RECT 121.660 14.365 122.335 14.525 ;
        RECT 119.150 14.165 119.810 14.195 ;
        RECT 119.150 13.945 119.985 14.165 ;
        RECT 119.640 13.865 119.985 13.945 ;
        RECT 118.810 13.585 119.465 13.755 ;
        RECT 118.810 12.955 119.045 13.415 ;
        RECT 119.215 13.215 119.465 13.585 ;
        RECT 119.815 13.335 119.985 13.865 ;
        RECT 120.155 13.905 120.695 14.275 ;
        RECT 121.030 14.185 121.435 14.355 ;
        RECT 120.155 13.505 120.395 13.905 ;
        RECT 120.875 13.735 121.095 14.015 ;
        RECT 120.565 13.565 121.095 13.735 ;
        RECT 120.565 13.335 120.735 13.565 ;
        RECT 121.265 13.405 121.435 14.185 ;
        RECT 121.605 13.575 121.955 14.195 ;
        RECT 122.125 13.575 122.335 14.365 ;
        RECT 122.525 14.395 124.025 14.565 ;
        RECT 122.525 13.705 122.695 14.395 ;
        RECT 124.385 14.225 124.555 15.005 ;
        RECT 125.360 14.875 125.530 15.005 ;
        RECT 122.865 14.055 124.555 14.225 ;
        RECT 124.725 14.445 125.190 14.835 ;
        RECT 125.360 14.705 125.755 14.875 ;
        RECT 122.865 13.875 123.035 14.055 ;
        RECT 119.815 13.165 120.735 13.335 ;
        RECT 120.905 12.955 121.095 13.395 ;
        RECT 121.265 13.125 122.215 13.405 ;
        RECT 122.525 13.315 122.785 13.705 ;
        RECT 123.205 13.635 123.995 13.885 ;
        RECT 122.435 13.145 122.785 13.315 ;
        RECT 122.995 12.955 123.325 13.415 ;
        RECT 124.200 13.345 124.370 14.055 ;
        RECT 124.725 13.855 124.895 14.445 ;
        RECT 124.540 13.635 124.895 13.855 ;
        RECT 125.065 13.635 125.415 14.255 ;
        RECT 125.585 13.345 125.755 14.705 ;
        RECT 126.120 14.535 126.445 15.320 ;
        RECT 125.925 13.485 126.385 14.535 ;
        RECT 124.200 13.175 125.055 13.345 ;
        RECT 125.260 13.175 125.755 13.345 ;
        RECT 125.925 12.955 126.255 13.315 ;
        RECT 126.615 13.215 126.785 15.335 ;
        RECT 126.955 15.005 127.285 15.505 ;
        RECT 127.455 14.835 127.710 15.335 ;
        RECT 126.960 14.665 127.710 14.835 ;
        RECT 126.960 13.675 127.190 14.665 ;
        RECT 127.360 14.490 127.710 14.495 ;
        RECT 130.570 14.490 131.400 14.500 ;
        RECT 127.360 13.850 131.400 14.490 ;
        RECT 127.360 13.845 127.710 13.850 ;
        RECT 130.570 13.820 131.400 13.850 ;
        RECT 126.960 13.505 127.710 13.675 ;
        RECT 126.955 12.955 127.285 13.335 ;
        RECT 127.455 13.215 127.710 13.505 ;
        RECT 116.760 12.785 127.800 12.955 ;
      LAYER mcon ;
        RECT 116.675 22.915 116.845 23.085 ;
        RECT 117.135 22.915 117.305 23.085 ;
        RECT 117.595 22.915 117.765 23.085 ;
        RECT 118.055 22.915 118.225 23.085 ;
        RECT 118.515 22.915 118.685 23.085 ;
        RECT 118.975 22.915 119.145 23.085 ;
        RECT 119.435 22.915 119.605 23.085 ;
        RECT 119.895 22.915 120.065 23.085 ;
        RECT 120.355 22.915 120.525 23.085 ;
        RECT 120.815 22.915 120.985 23.085 ;
        RECT 121.275 22.915 121.445 23.085 ;
        RECT 121.735 22.915 121.905 23.085 ;
        RECT 122.195 22.915 122.365 23.085 ;
        RECT 122.655 22.915 122.825 23.085 ;
        RECT 123.115 22.915 123.285 23.085 ;
        RECT 123.575 22.915 123.745 23.085 ;
        RECT 124.035 22.915 124.205 23.085 ;
        RECT 124.495 22.915 124.665 23.085 ;
        RECT 124.955 22.915 125.125 23.085 ;
        RECT 125.415 22.915 125.585 23.085 ;
        RECT 125.875 22.915 126.045 23.085 ;
        RECT 126.335 22.915 126.505 23.085 ;
        RECT 126.795 22.915 126.965 23.085 ;
        RECT 127.255 22.915 127.425 23.085 ;
        RECT 115.540 20.630 116.470 21.120 ;
        RECT 118.080 21.400 118.400 21.970 ;
        RECT 121.375 22.065 121.545 22.235 ;
        RECT 120.295 21.360 120.465 21.530 ;
        RECT 119.995 21.045 120.165 21.215 ;
        RECT 121.375 21.385 121.545 21.555 ;
        RECT 124.495 22.065 124.665 22.235 ;
        RECT 123.235 21.045 123.405 21.215 ;
        RECT 123.595 21.045 123.765 21.215 ;
        RECT 124.955 21.385 125.125 21.555 ;
        RECT 126.385 22.065 126.555 22.235 ;
        RECT 126.790 21.385 126.960 21.555 ;
        RECT 116.675 20.195 116.845 20.365 ;
        RECT 117.135 20.195 117.305 20.365 ;
        RECT 117.595 20.195 117.765 20.365 ;
        RECT 118.055 20.195 118.225 20.365 ;
        RECT 118.515 20.195 118.685 20.365 ;
        RECT 118.975 20.195 119.145 20.365 ;
        RECT 119.435 20.195 119.605 20.365 ;
        RECT 119.895 20.195 120.065 20.365 ;
        RECT 120.355 20.195 120.525 20.365 ;
        RECT 120.815 20.195 120.985 20.365 ;
        RECT 121.275 20.195 121.445 20.365 ;
        RECT 121.735 20.195 121.905 20.365 ;
        RECT 122.195 20.195 122.365 20.365 ;
        RECT 122.655 20.195 122.825 20.365 ;
        RECT 123.115 20.195 123.285 20.365 ;
        RECT 123.575 20.195 123.745 20.365 ;
        RECT 124.035 20.195 124.205 20.365 ;
        RECT 124.495 20.195 124.665 20.365 ;
        RECT 124.955 20.195 125.125 20.365 ;
        RECT 125.415 20.195 125.585 20.365 ;
        RECT 125.875 20.195 126.045 20.365 ;
        RECT 126.335 20.195 126.505 20.365 ;
        RECT 126.795 20.195 126.965 20.365 ;
        RECT 127.255 20.195 127.425 20.365 ;
        RECT 118.075 19.215 118.245 19.385 ;
        RECT 118.535 19.215 118.705 19.385 ;
        RECT 118.995 19.215 119.165 19.385 ;
        RECT 119.455 19.215 119.625 19.385 ;
        RECT 119.915 19.215 120.085 19.385 ;
        RECT 120.375 19.215 120.545 19.385 ;
        RECT 118.910 17.660 119.250 17.970 ;
        RECT 123.245 19.165 123.415 19.335 ;
        RECT 123.705 19.165 123.875 19.335 ;
        RECT 124.165 19.165 124.335 19.335 ;
        RECT 124.625 19.165 124.795 19.335 ;
        RECT 125.085 19.165 125.255 19.335 ;
        RECT 118.075 16.495 118.245 16.665 ;
        RECT 118.535 16.495 118.705 16.665 ;
        RECT 118.995 16.495 119.165 16.665 ;
        RECT 119.455 16.495 119.625 16.665 ;
        RECT 119.915 16.495 120.085 16.665 ;
        RECT 120.375 16.495 120.545 16.665 ;
        RECT 123.245 16.445 123.415 16.615 ;
        RECT 123.705 16.445 123.875 16.615 ;
        RECT 124.165 16.445 124.335 16.615 ;
        RECT 124.625 16.445 124.795 16.615 ;
        RECT 125.085 16.445 125.255 16.615 ;
        RECT 116.905 15.505 117.075 15.675 ;
        RECT 117.365 15.505 117.535 15.675 ;
        RECT 117.825 15.505 117.995 15.675 ;
        RECT 118.285 15.505 118.455 15.675 ;
        RECT 118.745 15.505 118.915 15.675 ;
        RECT 119.205 15.505 119.375 15.675 ;
        RECT 119.665 15.505 119.835 15.675 ;
        RECT 120.125 15.505 120.295 15.675 ;
        RECT 120.585 15.505 120.755 15.675 ;
        RECT 121.045 15.505 121.215 15.675 ;
        RECT 121.505 15.505 121.675 15.675 ;
        RECT 121.965 15.505 122.135 15.675 ;
        RECT 122.425 15.505 122.595 15.675 ;
        RECT 122.885 15.505 123.055 15.675 ;
        RECT 123.345 15.505 123.515 15.675 ;
        RECT 123.805 15.505 123.975 15.675 ;
        RECT 124.265 15.505 124.435 15.675 ;
        RECT 124.725 15.505 124.895 15.675 ;
        RECT 125.185 15.505 125.355 15.675 ;
        RECT 125.645 15.505 125.815 15.675 ;
        RECT 126.105 15.505 126.275 15.675 ;
        RECT 126.565 15.505 126.735 15.675 ;
        RECT 127.025 15.505 127.195 15.675 ;
        RECT 127.485 15.505 127.655 15.675 ;
        RECT 118.340 13.890 118.630 14.530 ;
        RECT 121.605 14.655 121.775 14.825 ;
        RECT 120.525 13.950 120.695 14.120 ;
        RECT 120.225 13.635 120.395 13.805 ;
        RECT 121.605 13.975 121.775 14.145 ;
        RECT 124.725 14.655 124.895 14.825 ;
        RECT 123.465 13.635 123.635 13.805 ;
        RECT 123.825 13.635 123.995 13.805 ;
        RECT 125.185 13.975 125.355 14.145 ;
        RECT 126.615 14.655 126.785 14.825 ;
        RECT 127.020 13.975 127.190 14.145 ;
        RECT 116.905 12.785 117.075 12.955 ;
        RECT 117.365 12.785 117.535 12.955 ;
        RECT 117.825 12.785 117.995 12.955 ;
        RECT 118.285 12.785 118.455 12.955 ;
        RECT 118.745 12.785 118.915 12.955 ;
        RECT 119.205 12.785 119.375 12.955 ;
        RECT 119.665 12.785 119.835 12.955 ;
        RECT 120.125 12.785 120.295 12.955 ;
        RECT 120.585 12.785 120.755 12.955 ;
        RECT 121.045 12.785 121.215 12.955 ;
        RECT 121.505 12.785 121.675 12.955 ;
        RECT 121.965 12.785 122.135 12.955 ;
        RECT 122.425 12.785 122.595 12.955 ;
        RECT 122.885 12.785 123.055 12.955 ;
        RECT 123.345 12.785 123.515 12.955 ;
        RECT 123.805 12.785 123.975 12.955 ;
        RECT 124.265 12.785 124.435 12.955 ;
        RECT 124.725 12.785 124.895 12.955 ;
        RECT 125.185 12.785 125.355 12.955 ;
        RECT 125.645 12.785 125.815 12.955 ;
        RECT 126.105 12.785 126.275 12.955 ;
        RECT 126.565 12.785 126.735 12.955 ;
        RECT 127.025 12.785 127.195 12.955 ;
        RECT 127.485 12.785 127.655 12.955 ;
      LAYER met1 ;
        RECT 0.590 24.295 3.050 25.730 ;
        RECT 128.090 24.295 129.300 24.400 ;
        RECT 0.590 23.085 129.300 24.295 ;
        RECT 0.590 20.810 3.050 23.085 ;
        RECT 116.530 22.760 129.300 23.085 ;
        RECT 121.315 22.220 121.605 22.265 ;
        RECT 124.435 22.220 124.725 22.265 ;
        RECT 126.325 22.220 126.615 22.265 ;
        RECT 110.500 22.020 114.690 22.170 ;
        RECT 121.315 22.080 126.615 22.220 ;
        RECT 121.315 22.035 121.605 22.080 ;
        RECT 124.435 22.035 124.725 22.080 ;
        RECT 126.325 22.035 126.615 22.080 ;
        RECT 118.050 22.020 118.430 22.030 ;
        RECT 110.500 21.380 118.430 22.020 ;
        RECT 110.500 21.170 114.690 21.380 ;
        RECT 118.050 21.340 118.430 21.380 ;
        RECT 120.235 21.245 120.525 21.560 ;
        RECT 121.315 21.540 121.605 21.585 ;
        RECT 124.895 21.540 125.185 21.585 ;
        RECT 126.730 21.540 127.020 21.585 ;
        RECT 121.315 21.400 127.020 21.540 ;
        RECT 121.315 21.355 121.605 21.400 ;
        RECT 124.895 21.355 125.185 21.400 ;
        RECT 126.730 21.355 127.020 21.400 ;
        RECT 119.935 21.200 120.525 21.245 ;
        RECT 122.295 21.200 122.855 21.220 ;
        RECT 123.175 21.200 123.825 21.245 ;
        RECT 110.500 3.180 111.500 21.170 ;
        RECT 113.780 18.530 114.580 21.170 ;
        RECT 115.130 20.530 116.670 21.150 ;
        RECT 119.935 21.060 123.825 21.200 ;
        RECT 119.935 21.015 120.225 21.060 ;
        RECT 122.295 20.890 122.855 21.060 ;
        RECT 123.175 21.015 123.825 21.060 ;
        RECT 115.120 20.520 116.740 20.530 ;
        RECT 115.120 20.040 127.570 20.520 ;
        RECT 113.460 17.580 114.630 18.530 ;
        RECT 115.120 17.600 116.450 20.040 ;
        RECT 128.090 19.660 129.300 22.760 ;
        RECT 130.480 22.060 131.480 22.130 ;
        RECT 130.480 21.910 157.390 22.060 ;
        RECT 130.190 21.240 157.390 21.910 ;
        RECT 130.480 21.130 157.390 21.240 ;
        RECT 130.810 21.000 157.390 21.130 ;
        RECT 120.510 19.540 123.310 19.560 ;
        RECT 117.930 19.490 123.310 19.540 ;
        RECT 124.330 19.490 125.420 19.500 ;
        RECT 128.090 19.490 129.350 19.660 ;
        RECT 117.930 19.060 129.350 19.490 ;
        RECT 120.510 19.020 129.350 19.060 ;
        RECT 123.100 19.010 129.350 19.020 ;
        RECT 125.370 18.990 129.350 19.010 ;
        RECT 128.090 18.920 129.350 18.990 ;
        RECT 118.850 17.920 119.310 18.000 ;
        RECT 118.850 17.630 119.350 17.920 ;
        RECT 115.120 17.570 116.910 17.600 ;
        RECT 118.910 17.580 119.350 17.630 ;
        RECT 120.820 17.870 121.780 17.940 ;
        RECT 120.820 17.590 121.790 17.870 ;
        RECT 115.120 16.820 117.990 17.570 ;
        RECT 120.820 17.560 121.780 17.590 ;
        RECT 125.640 17.380 126.490 18.110 ;
        RECT 119.925 16.820 120.295 16.830 ;
        RECT 115.120 16.770 123.190 16.820 ;
        RECT 115.120 16.290 125.400 16.770 ;
        RECT 115.120 16.280 123.190 16.290 ;
        RECT 113.170 14.680 114.480 15.140 ;
        RECT 113.170 14.600 114.490 14.680 ;
        RECT 113.170 13.850 114.890 14.600 ;
        RECT 113.170 13.630 114.480 13.850 ;
        RECT 115.120 13.810 116.450 16.280 ;
        RECT 116.760 15.830 116.910 15.850 ;
        RECT 128.090 15.830 129.300 18.920 ;
        RECT 116.760 15.360 129.300 15.830 ;
        RECT 116.760 15.350 127.800 15.360 ;
        RECT 128.090 15.320 129.300 15.360 ;
        RECT 121.545 14.810 121.835 14.855 ;
        RECT 124.665 14.810 124.955 14.855 ;
        RECT 126.555 14.810 126.845 14.855 ;
        RECT 121.545 14.670 126.845 14.810 ;
        RECT 121.545 14.625 121.835 14.670 ;
        RECT 124.665 14.625 124.955 14.670 ;
        RECT 126.555 14.625 126.845 14.670 ;
        RECT 130.680 14.625 131.680 14.710 ;
        RECT 118.310 14.530 118.660 14.590 ;
        RECT 130.680 14.530 135.175 14.625 ;
        RECT 116.630 13.900 118.660 14.530 ;
        RECT 118.310 13.830 118.660 13.900 ;
        RECT 120.465 13.835 120.755 14.150 ;
        RECT 121.545 14.130 121.835 14.175 ;
        RECT 125.125 14.130 125.415 14.175 ;
        RECT 126.960 14.130 127.250 14.175 ;
        RECT 121.545 13.990 127.250 14.130 ;
        RECT 121.545 13.945 121.835 13.990 ;
        RECT 125.125 13.945 125.415 13.990 ;
        RECT 126.960 13.945 127.250 13.990 ;
        RECT 115.120 13.120 116.490 13.810 ;
        RECT 120.165 13.790 120.755 13.835 ;
        RECT 121.900 13.790 122.450 13.800 ;
        RECT 123.405 13.790 124.055 13.835 ;
        RECT 130.510 13.790 135.175 14.530 ;
        RECT 120.165 13.650 124.055 13.790 ;
        RECT 130.680 13.710 135.175 13.790 ;
        RECT 131.075 13.695 135.175 13.710 ;
        RECT 120.165 13.605 120.455 13.650 ;
        RECT 121.900 13.530 122.450 13.650 ;
        RECT 123.405 13.605 124.055 13.650 ;
        RECT 115.120 13.110 116.820 13.120 ;
        RECT 115.120 12.630 127.800 13.110 ;
        RECT 115.120 11.710 116.450 12.630 ;
        RECT 114.980 10.030 116.580 11.710 ;
        RECT 134.245 4.795 135.175 13.695 ;
        RECT 134.245 3.550 135.180 4.795 ;
        RECT 111.890 3.180 113.270 3.350 ;
        RECT 110.500 2.250 113.270 3.180 ;
        RECT 111.500 2.180 113.270 2.250 ;
        RECT 111.890 2.140 113.270 2.180 ;
        RECT 134.020 1.370 135.480 3.550 ;
        RECT 156.330 3.540 157.390 21.000 ;
        RECT 156.080 1.790 157.610 3.540 ;
        RECT 134.245 1.295 135.180 1.370 ;
        RECT 134.245 1.255 135.175 1.295 ;
      LAYER via ;
        RECT 0.640 20.810 3.000 25.730 ;
        RECT 122.345 20.890 122.805 21.220 ;
        RECT 124.380 19.010 125.370 19.500 ;
        RECT 128.160 18.920 129.300 19.660 ;
        RECT 118.960 17.580 119.300 17.920 ;
        RECT 125.700 17.410 126.430 18.080 ;
        RECT 113.220 13.630 114.430 15.140 ;
        RECT 114.470 13.850 114.840 14.600 ;
        RECT 116.690 13.900 117.150 14.520 ;
        RECT 121.950 13.530 122.400 13.800 ;
        RECT 115.030 10.030 116.530 11.710 ;
        RECT 111.940 2.140 113.220 3.350 ;
        RECT 134.070 1.370 135.430 3.550 ;
        RECT 156.130 1.790 157.560 3.540 ;
      LAYER met2 ;
        RECT 0.640 20.760 3.000 25.780 ;
        RECT 122.345 21.220 122.805 21.270 ;
        RECT 122.345 20.840 122.815 21.220 ;
        RECT 122.355 20.040 122.815 20.840 ;
        RECT 125.720 20.040 126.430 20.050 ;
        RECT 122.350 19.700 126.430 20.040 ;
        RECT 124.380 18.960 125.370 19.550 ;
        RECT 125.720 18.290 126.430 19.700 ;
        RECT 128.160 18.870 129.300 19.710 ;
        RECT 125.720 18.130 126.440 18.290 ;
        RECT 118.960 17.910 119.300 17.970 ;
        RECT 118.950 16.130 119.330 17.910 ;
        RECT 125.700 17.360 126.440 18.130 ;
        RECT 125.760 16.190 126.440 17.360 ;
        RECT 116.720 15.900 119.330 16.130 ;
        RECT 90.130 14.820 91.260 15.530 ;
        RECT 113.220 14.820 114.430 15.190 ;
        RECT 90.130 13.820 114.430 14.820 ;
        RECT 90.130 13.650 91.260 13.820 ;
        RECT 113.220 13.580 114.430 13.820 ;
        RECT 114.470 14.550 114.840 14.650 ;
        RECT 116.720 14.570 117.120 15.900 ;
        RECT 121.950 15.860 126.450 16.190 ;
        RECT 116.690 14.550 117.150 14.570 ;
        RECT 114.470 13.880 117.150 14.550 ;
        RECT 114.470 13.800 114.840 13.880 ;
        RECT 116.690 13.850 117.150 13.880 ;
        RECT 121.950 13.850 122.390 15.860 ;
        RECT 121.950 13.480 122.400 13.850 ;
        RECT 115.030 9.980 116.530 11.760 ;
        RECT 111.940 2.090 113.220 3.400 ;
        RECT 134.070 1.320 135.430 3.600 ;
        RECT 156.130 1.740 157.560 3.590 ;
      LAYER via2 ;
        RECT 0.640 20.810 3.000 25.730 ;
        RECT 90.130 13.700 91.260 15.480 ;
        RECT 115.030 10.030 116.530 11.710 ;
        RECT 111.940 2.140 113.220 3.350 ;
        RECT 134.070 1.370 135.430 3.550 ;
        RECT 156.130 1.790 157.560 3.540 ;
      LAYER met3 ;
        RECT 0.590 20.785 3.050 25.755 ;
        RECT 90.080 13.675 91.310 15.505 ;
        RECT 86.880 10.110 100.230 11.610 ;
        RECT 114.980 10.005 116.580 11.735 ;
        RECT 111.890 2.115 113.270 3.375 ;
        RECT 134.020 1.345 135.480 3.575 ;
        RECT 156.080 1.765 157.610 3.565 ;
      LAYER via3 ;
        RECT 0.640 20.810 3.000 25.730 ;
        RECT 90.130 13.700 91.260 15.480 ;
        RECT 86.885 10.115 88.375 11.605 ;
        RECT 98.700 10.110 100.200 11.610 ;
        RECT 115.030 10.030 116.530 11.710 ;
        RECT 111.940 2.140 113.220 3.350 ;
        RECT 134.070 1.370 135.430 3.550 ;
        RECT 156.130 1.790 157.560 3.540 ;
      LAYER met4 ;
        RECT 0.635 20.805 1.000 25.735 ;
        RECT 2.500 20.805 3.005 25.735 ;
        RECT 90.125 13.695 91.265 15.485 ;
        RECT 50.500 10.110 88.380 11.610 ;
        RECT 90.320 1.000 90.920 13.695 ;
        RECT 98.695 11.610 100.205 11.615 ;
        RECT 115.025 11.610 116.535 11.715 ;
        RECT 98.695 10.110 116.535 11.610 ;
        RECT 98.695 10.105 100.205 10.110 ;
        RECT 115.025 10.025 116.535 10.110 ;
        RECT 111.935 2.135 113.225 3.355 ;
        RECT 112.400 1.000 113.000 2.135 ;
        RECT 134.065 1.365 135.435 3.555 ;
        RECT 156.125 1.785 157.565 3.545 ;
        RECT 134.480 1.000 135.080 1.365 ;
        RECT 156.560 1.000 157.160 1.785 ;
  END
END tt_um_vks_pll
END LIBRARY

