VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_vks_pll
  CLASS BLOCK ;
  FOREIGN tt_um_vks_pll ;
  ORIGIN 0.000 0.000 ;
  SIZE 161.000 BY 225.760 ;
  PIN clk
    PORT
      LAYER met4 ;
        RECT 154.870 224.760 155.170 225.760 ;
    END
  END clk
  PIN ena
    PORT
      LAYER met4 ;
        RECT 158.550 224.760 158.850 225.760 ;
    END
  END ena
  PIN rst_n
    PORT
      LAYER met4 ;
        RECT 151.190 224.760 151.490 225.760 ;
    END
  END rst_n
  PIN ua[0]
    ANTENNAGATEAREA 5.400000 ;
    PORT
      LAYER met4 ;
        RECT 156.560 0.000 157.160 1.000 ;
    END
  END ua[0]
  PIN ua[1]
    ANTENNADIFFAREA 0.580000 ;
    PORT
      LAYER met4 ;
        RECT 134.480 0.000 135.080 1.000 ;
    END
  END ua[1]
  PIN ua[2]
    ANTENNAGATEAREA 20.799999 ;
    PORT
      LAYER met4 ;
        RECT 112.400 0.000 113.000 1.000 ;
    END
  END ua[2]
  PIN ua[3]
    ANTENNADIFFAREA 2.022500 ;
    PORT
      LAYER met4 ;
        RECT 90.320 0.000 90.920 1.000 ;
    END
  END ua[3]
  PIN ua[4]
    ANTENNAGATEAREA 0.300000 ;
    PORT
      LAYER met4 ;
        RECT 68.240 0.000 68.840 1.000 ;
    END
  END ua[4]
  PIN ua[5]
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 46.160 0.000 46.760 1.000 ;
    END
  END ua[5]
  PIN ua[6]
    PORT
      LAYER met4 ;
        RECT 24.080 0.000 24.680 1.000 ;
    END
  END ua[6]
  PIN ua[7]
    PORT
      LAYER met4 ;
        RECT 2.000 0.000 2.600 1.000 ;
    END
  END ua[7]
  PIN ui_in[0]
    ANTENNAGATEAREA 2.000000 ;
    PORT
      LAYER met4 ;
        RECT 147.510 224.750 147.810 225.750 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    ANTENNAGATEAREA 5.000000 ;
    PORT
      LAYER met4 ;
        RECT 143.830 224.760 144.130 225.760 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met4 ;
        RECT 140.150 224.760 140.450 225.760 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met4 ;
        RECT 136.470 224.760 136.770 225.760 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met4 ;
        RECT 132.790 224.760 133.090 225.760 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    PORT
      LAYER met4 ;
        RECT 129.110 224.760 129.410 225.760 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met4 ;
        RECT 125.430 224.760 125.730 225.760 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    PORT
      LAYER met4 ;
        RECT 121.750 224.760 122.050 225.760 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met4 ;
        RECT 118.070 224.760 118.370 225.760 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    PORT
      LAYER met4 ;
        RECT 114.390 224.760 114.690 225.760 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met4 ;
        RECT 110.710 224.760 111.010 225.760 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met4 ;
        RECT 107.030 224.760 107.330 225.760 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    PORT
      LAYER met4 ;
        RECT 103.350 224.760 103.650 225.760 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    PORT
      LAYER met4 ;
        RECT 99.670 224.760 99.970 225.760 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met4 ;
        RECT 95.990 224.760 96.290 225.760 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met4 ;
        RECT 92.310 224.760 92.610 225.760 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    ANTENNADIFFAREA 104.138847 ;
    PORT
      LAYER met4 ;
        RECT 29.750 224.760 30.050 225.760 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    ANTENNAGATEAREA 0.756000 ;
    ANTENNADIFFAREA 133.305695 ;
    PORT
      LAYER met4 ;
        RECT 26.070 224.760 26.370 225.760 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    ANTENNADIFFAREA 104.138847 ;
    PORT
      LAYER met4 ;
        RECT 22.390 224.760 22.690 225.760 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    ANTENNADIFFAREA 104.138847 ;
    PORT
      LAYER met4 ;
        RECT 18.710 224.760 19.010 225.760 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    ANTENNAGATEAREA 0.756000 ;
    ANTENNADIFFAREA 133.305695 ;
    PORT
      LAYER met4 ;
        RECT 15.030 224.760 15.330 225.760 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    ANTENNAGATEAREA 0.756000 ;
    ANTENNADIFFAREA 133.305695 ;
    PORT
      LAYER met4 ;
        RECT 11.350 224.760 11.650 225.760 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    ANTENNADIFFAREA 104.138847 ;
    PORT
      LAYER met4 ;
        RECT 7.670 224.760 7.970 225.760 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    ANTENNADIFFAREA 104.138847 ;
    PORT
      LAYER met4 ;
        RECT 3.990 224.760 4.290 225.760 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    PORT
      LAYER met4 ;
        RECT 59.190 224.760 59.490 225.760 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 55.510 224.760 55.810 225.760 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    PORT
      LAYER met4 ;
        RECT 51.830 224.760 52.130 225.760 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    PORT
      LAYER met4 ;
        RECT 48.150 224.760 48.450 225.760 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met4 ;
        RECT 44.470 224.760 44.770 225.760 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met4 ;
        RECT 40.790 224.760 41.090 225.760 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    PORT
      LAYER met4 ;
        RECT 37.110 224.760 37.410 225.760 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    PORT
      LAYER met4 ;
        RECT 33.430 224.760 33.730 225.760 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.511500 ;
    PORT
      LAYER met4 ;
        RECT 88.630 224.760 88.930 225.760 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.511500 ;
    PORT
      LAYER met4 ;
        RECT 84.950 224.760 85.250 225.760 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 81.270 224.760 81.570 225.760 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 77.590 224.760 77.890 225.760 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    PORT
      LAYER met4 ;
        RECT 73.910 224.760 74.210 225.760 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    PORT
      LAYER met4 ;
        RECT 70.230 224.760 70.530 225.760 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    PORT
      LAYER met4 ;
        RECT 66.550 224.760 66.850 225.760 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    PORT
      LAYER met4 ;
        RECT 62.870 224.760 63.170 225.760 ;
    END
  END uo_out[7]
  PIN VPWR
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1.000 5.000 2.500 220.760 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 49.000 5.000 50.500 220.760 ;
    END
  END VGND
  OBS
      LAYER nwell ;
        RECT 56.330 220.700 57.570 220.710 ;
        RECT 56.330 219.260 77.490 220.700 ;
        RECT 57.570 219.095 77.490 219.260 ;
        RECT 133.180 219.590 134.720 220.270 ;
      LAYER pwell ;
        RECT 56.940 217.870 57.620 218.860 ;
        RECT 57.815 217.895 60.005 218.805 ;
        RECT 60.495 217.895 62.685 218.805 ;
        RECT 63.175 217.895 65.365 218.805 ;
        RECT 65.910 218.575 68.190 218.805 ;
        RECT 71.395 218.575 72.325 218.795 ;
        RECT 65.910 217.895 76.835 218.575 ;
        RECT 76.855 217.980 77.285 218.765 ;
        RECT 59.745 217.705 59.915 217.895 ;
        RECT 62.425 217.705 62.595 217.895 ;
        RECT 65.105 217.705 65.275 217.895 ;
        RECT 76.525 217.705 76.695 217.895 ;
      LAYER nwell ;
        RECT 62.150 215.910 69.210 217.360 ;
        RECT 63.390 215.755 69.210 215.910 ;
      LAYER pwell ;
        RECT 63.060 214.535 63.740 215.430 ;
        RECT 64.735 215.375 66.325 215.465 ;
        RECT 63.755 214.555 66.325 215.375 ;
        RECT 66.775 214.555 68.965 215.465 ;
        RECT 63.755 214.535 63.895 214.555 ;
        RECT 63.060 214.440 63.895 214.535 ;
        RECT 63.725 214.365 63.895 214.440 ;
        RECT 66.865 214.365 67.035 214.555 ;
        RECT 10.565 213.835 10.735 214.025 ;
        RECT 23.365 213.845 23.535 214.035 ;
        RECT 35.275 213.845 35.445 214.035 ;
        RECT 10.425 213.155 19.155 213.835 ;
        RECT 13.940 212.935 14.850 213.155 ;
        RECT 16.390 212.925 19.155 213.155 ;
        RECT 19.170 212.880 20.080 213.770 ;
        RECT 23.225 213.165 31.955 213.845 ;
        RECT 26.740 212.945 27.650 213.165 ;
        RECT 29.190 212.935 31.955 213.165 ;
        RECT 31.980 212.820 32.890 213.710 ;
        RECT 35.135 213.165 43.865 213.845 ;
        RECT 38.650 212.945 39.560 213.165 ;
        RECT 41.100 212.935 43.865 213.165 ;
        RECT 43.880 212.850 44.790 213.740 ;
      LAYER nwell ;
        RECT 10.230 212.580 19.350 212.635 ;
        RECT 10.230 211.510 20.430 212.580 ;
        RECT 23.030 212.540 32.150 212.645 ;
        RECT 10.230 211.030 19.350 211.510 ;
        RECT 23.030 211.500 33.440 212.540 ;
        RECT 34.940 212.000 44.060 212.645 ;
        RECT 59.200 212.570 77.490 214.020 ;
        RECT 60.440 212.415 77.490 212.570 ;
        RECT 23.030 211.040 32.150 211.500 ;
        RECT 34.940 211.040 44.940 212.000 ;
      LAYER pwell ;
        RECT 59.770 211.190 60.450 212.180 ;
        RECT 60.685 211.215 62.875 212.125 ;
        RECT 63.365 211.215 65.555 212.125 ;
        RECT 65.910 211.895 68.190 212.125 ;
        RECT 71.395 211.895 72.325 212.115 ;
        RECT 65.910 211.215 76.835 211.895 ;
        RECT 76.855 211.300 77.285 212.085 ;
      LAYER nwell ;
        RECT 43.900 210.890 44.940 211.040 ;
      LAYER pwell ;
        RECT 62.615 211.025 62.785 211.215 ;
        RECT 65.295 211.025 65.465 211.215 ;
        RECT 76.525 211.025 76.695 211.215 ;
      LAYER nwell ;
        RECT 85.280 206.100 86.400 206.420 ;
        RECT 85.280 204.890 117.670 206.100 ;
        RECT 86.400 204.495 117.670 204.890 ;
      LAYER pwell ;
        RECT 85.520 203.210 86.270 204.260 ;
        RECT 86.605 203.295 87.955 204.205 ;
        RECT 88.175 203.295 89.525 204.205 ;
        RECT 89.775 203.975 92.540 204.205 ;
        RECT 94.080 203.975 94.990 204.195 ;
        RECT 89.775 203.295 98.505 203.975 ;
        RECT 98.715 203.380 99.145 204.165 ;
        RECT 99.375 203.975 102.140 204.205 ;
        RECT 103.680 203.975 104.590 204.195 ;
        RECT 108.285 203.975 111.050 204.205 ;
        RECT 112.590 203.975 113.500 204.195 ;
        RECT 99.375 203.295 108.105 203.975 ;
        RECT 108.285 203.295 117.015 203.975 ;
        RECT 117.035 203.380 117.465 204.165 ;
        RECT 87.655 203.105 87.825 203.295 ;
        RECT 89.225 203.105 89.395 203.295 ;
        RECT 98.195 203.105 98.365 203.295 ;
        RECT 107.795 203.105 107.965 203.295 ;
        RECT 116.705 203.105 116.875 203.295 ;
      LAYER nwell ;
        RECT 10.950 201.730 21.590 202.570 ;
        RECT 23.370 202.560 33.410 202.570 ;
        RECT 10.950 200.965 20.990 201.730 ;
        RECT 23.370 201.220 34.370 202.560 ;
        RECT 45.720 202.550 47.100 202.560 ;
        RECT 23.370 200.965 33.410 201.220 ;
        RECT 35.690 200.960 47.100 202.550 ;
        RECT 35.690 200.945 45.730 200.960 ;
      LAYER pwell ;
        RECT 14.660 200.445 15.570 200.665 ;
        RECT 17.110 200.445 20.795 200.675 ;
        RECT 11.145 199.765 20.795 200.445 ;
        RECT 20.890 199.870 21.500 200.720 ;
        RECT 27.080 200.445 27.990 200.665 ;
        RECT 29.530 200.445 33.215 200.675 ;
        RECT 23.565 199.765 33.215 200.445 ;
        RECT 33.530 199.840 34.290 200.560 ;
        RECT 39.400 200.425 40.310 200.645 ;
        RECT 41.850 200.425 45.535 200.655 ;
        RECT 11.285 199.575 11.455 199.765 ;
        RECT 23.705 199.575 23.875 199.765 ;
        RECT 35.885 199.745 45.535 200.425 ;
        RECT 36.025 199.555 36.195 199.745 ;
        RECT 45.600 199.730 46.390 200.610 ;
      LAYER nwell ;
        RECT 95.710 196.650 97.250 196.690 ;
        RECT 95.710 195.045 108.260 196.650 ;
        RECT 95.710 195.000 97.250 195.045 ;
      LAYER pwell ;
        RECT 96.280 193.790 97.060 194.750 ;
        RECT 97.140 194.525 99.420 194.755 ;
        RECT 102.625 194.525 103.555 194.745 ;
        RECT 97.140 193.845 108.065 194.525 ;
        RECT 107.755 193.655 107.925 193.845 ;
      LAYER nwell ;
        RECT 97.860 192.300 98.770 192.310 ;
        RECT 97.860 192.280 103.320 192.300 ;
        RECT 97.860 191.320 105.880 192.280 ;
        RECT 98.580 190.695 105.880 191.320 ;
        RECT 101.540 190.680 105.880 190.695 ;
        RECT 103.200 190.675 105.880 190.680 ;
      LAYER pwell ;
        RECT 98.070 189.490 98.930 190.450 ;
        RECT 99.925 190.315 101.515 190.405 ;
        RECT 98.945 189.495 101.515 190.315 ;
        RECT 98.945 189.475 99.085 189.495 ;
        RECT 103.445 189.475 105.635 190.385 ;
        RECT 98.915 189.305 99.085 189.475 ;
        RECT 103.535 189.285 103.705 189.475 ;
      LAYER nwell ;
        RECT 133.180 189.320 134.785 219.590 ;
      LAYER pwell ;
        RECT 135.075 215.710 135.985 219.395 ;
        RECT 135.305 214.170 135.985 215.710 ;
        RECT 135.085 213.260 135.985 214.170 ;
        RECT 135.305 210.055 135.985 213.260 ;
        RECT 135.305 209.885 136.175 210.055 ;
        RECT 135.305 209.745 135.985 209.885 ;
        RECT 135.115 209.295 135.900 209.725 ;
        RECT 135.075 205.590 135.985 209.275 ;
        RECT 135.305 204.050 135.985 205.590 ;
        RECT 135.085 203.140 135.985 204.050 ;
        RECT 135.305 199.935 135.985 203.140 ;
        RECT 135.305 199.765 136.175 199.935 ;
        RECT 135.305 199.625 135.985 199.765 ;
        RECT 135.115 199.175 135.900 199.605 ;
        RECT 135.075 195.480 135.985 199.165 ;
        RECT 135.305 193.940 135.985 195.480 ;
        RECT 135.085 193.030 135.985 193.940 ;
        RECT 135.305 189.825 135.985 193.030 ;
        RECT 135.305 189.655 136.175 189.825 ;
        RECT 135.305 189.515 135.985 189.655 ;
        RECT 135.260 189.430 136.050 189.480 ;
        RECT 135.250 188.700 136.050 189.430 ;
      LAYER nwell ;
        RECT 95.930 187.900 97.020 187.970 ;
        RECT 95.930 186.295 108.140 187.900 ;
        RECT 95.930 186.240 97.020 186.295 ;
      LAYER pwell ;
        RECT 96.180 185.100 96.860 185.930 ;
        RECT 97.020 185.775 99.300 186.005 ;
        RECT 102.505 185.775 103.435 185.995 ;
        RECT 97.020 185.095 107.945 185.775 ;
        RECT 107.635 184.905 107.805 185.095 ;
      LAYER nwell ;
        RECT 88.400 150.450 90.510 150.460 ;
        RECT 92.620 150.450 94.730 150.460 ;
        RECT 69.220 150.120 70.240 150.170 ;
        RECT 69.060 150.080 70.240 150.120 ;
        RECT 57.900 148.475 70.240 150.080 ;
        RECT 72.570 148.475 75.710 150.080 ;
        RECT 69.220 148.470 70.240 148.475 ;
      LAYER pwell ;
        RECT 62.605 147.955 63.535 148.175 ;
        RECT 66.740 147.955 69.020 148.185 ;
        RECT 58.095 147.275 69.020 147.955 ;
        RECT 69.040 147.380 70.300 148.290 ;
        RECT 72.815 147.275 75.005 148.185 ;
        RECT 75.075 147.360 75.505 148.145 ;
        RECT 58.235 147.085 58.405 147.275 ;
        RECT 72.905 147.085 73.075 147.275 ;
      LAYER nwell ;
        RECT 62.580 146.380 64.860 146.390 ;
        RECT 67.830 146.380 68.860 146.400 ;
        RECT 62.580 146.330 68.860 146.380 ;
        RECT 60.070 144.775 68.860 146.330 ;
        RECT 78.400 146.000 85.250 150.190 ;
        RECT 88.400 147.470 94.730 150.450 ;
        RECT 96.050 147.470 98.160 150.460 ;
      LAYER pwell ;
        RECT 98.240 147.530 102.100 150.330 ;
      LAYER nwell ;
        RECT 60.070 144.740 64.860 144.775 ;
        RECT 67.830 144.770 68.860 144.775 ;
        RECT 60.070 144.725 62.750 144.740 ;
      LAYER pwell ;
        RECT 60.315 143.525 62.505 144.435 ;
        RECT 64.985 144.395 66.575 144.485 ;
        RECT 64.985 143.575 67.555 144.395 ;
        RECT 67.740 143.710 68.870 144.450 ;
        RECT 67.415 143.555 67.555 143.575 ;
        RECT 62.245 143.335 62.415 143.525 ;
        RECT 67.415 143.385 67.585 143.555 ;
        RECT 78.450 142.820 85.800 145.820 ;
      LAYER nwell ;
        RECT 87.770 145.360 99.960 147.470 ;
      LAYER pwell ;
        RECT 92.920 143.990 99.920 145.310 ;
        RECT 100.020 143.990 103.880 146.090 ;
        RECT 92.920 143.760 103.880 143.990 ;
        RECT 92.920 143.300 99.920 143.760 ;
        RECT 100.020 143.290 103.880 143.760 ;
      LAYER nwell ;
        RECT 57.670 141.080 69.990 142.670 ;
        RECT 87.760 141.120 99.950 143.230 ;
        RECT 57.670 141.065 69.090 141.080 ;
      LAYER pwell ;
        RECT 62.375 140.545 63.305 140.765 ;
        RECT 66.510 140.545 68.790 140.775 ;
        RECT 57.865 139.865 68.790 140.545 ;
        RECT 58.005 139.675 58.175 139.865 ;
        RECT 69.090 139.620 70.000 140.990 ;
        RECT 92.900 139.740 99.900 141.060 ;
        RECT 100.000 139.740 103.860 141.850 ;
        RECT 92.900 139.430 103.860 139.740 ;
        RECT 92.900 139.050 99.900 139.430 ;
        RECT 100.000 139.050 103.860 139.430 ;
      LAYER nwell ;
        RECT 71.240 138.705 81.280 138.710 ;
        RECT 70.220 137.215 81.280 138.705 ;
        RECT 71.240 137.105 81.280 137.215 ;
      LAYER pwell ;
        RECT 70.790 135.820 71.420 136.900 ;
      LAYER nwell ;
        RECT 87.760 136.890 99.950 139.000 ;
        RECT 89.770 136.870 91.380 136.890 ;
      LAYER pwell ;
        RECT 71.435 136.585 75.120 136.815 ;
        RECT 76.660 136.585 77.570 136.805 ;
        RECT 71.435 135.905 81.085 136.585 ;
        RECT 80.775 135.715 80.945 135.905 ;
      LAYER nwell ;
        RECT 69.685 134.420 81.260 135.190 ;
        RECT 89.770 135.120 91.375 136.870 ;
      LAYER pwell ;
        RECT 91.665 136.545 92.575 136.675 ;
        RECT 91.665 136.375 92.765 136.545 ;
        RECT 91.665 135.325 92.575 136.375 ;
        RECT 92.910 134.820 99.910 136.830 ;
        RECT 100.010 134.810 103.870 137.610 ;
      LAYER nwell ;
        RECT 69.680 133.585 81.260 134.420 ;
        RECT 69.680 133.580 71.230 133.585 ;
      LAYER pwell ;
        RECT 70.790 132.310 71.400 133.420 ;
        RECT 71.415 133.065 75.100 133.295 ;
        RECT 76.640 133.065 77.550 133.285 ;
        RECT 71.415 132.385 81.065 133.065 ;
        RECT 80.755 132.195 80.925 132.385 ;
      LAYER nwell ;
        RECT 69.835 130.190 81.320 131.680 ;
        RECT 70.840 130.180 81.320 130.190 ;
        RECT 71.280 130.075 81.320 130.180 ;
      LAYER pwell ;
        RECT 70.800 128.740 71.390 129.940 ;
        RECT 71.475 129.555 75.160 129.785 ;
        RECT 76.700 129.555 77.610 129.775 ;
        RECT 71.475 128.875 81.125 129.555 ;
        RECT 84.570 128.950 111.810 132.020 ;
        RECT 80.815 128.685 80.985 128.875 ;
      LAYER nwell ;
        RECT 106.070 23.170 109.920 28.610 ;
        RECT 111.190 23.170 115.040 28.610 ;
        RECT 116.310 23.160 120.160 28.600 ;
        RECT 121.430 23.160 125.280 28.600 ;
        RECT 99.220 17.770 102.330 21.960 ;
        RECT 103.610 17.710 108.400 21.900 ;
        RECT 109.670 17.710 114.460 21.900 ;
        RECT 115.730 17.700 120.520 21.890 ;
      LAYER pwell ;
        RECT 121.440 17.240 125.190 22.490 ;
      LAYER nwell ;
        RECT 138.850 19.580 142.290 27.770 ;
        RECT 144.600 19.260 146.860 27.450 ;
        RECT 150.880 18.810 153.730 28.000 ;
      LAYER pwell ;
        RECT 99.640 12.870 102.170 17.120 ;
        RECT 104.440 12.940 108.090 17.190 ;
        RECT 110.530 12.920 114.180 17.170 ;
        RECT 116.540 12.930 120.190 17.180 ;
        RECT 137.115 14.065 139.275 18.065 ;
        RECT 140.865 14.525 143.025 18.525 ;
        RECT 144.150 13.860 146.510 16.560 ;
      LAYER nwell ;
        RECT 150.285 14.340 154.245 17.530 ;
      LAYER pwell ;
        RECT 104.400 7.080 108.150 12.330 ;
        RECT 110.500 7.080 114.250 12.330 ;
        RECT 116.580 7.100 120.330 12.350 ;
        RECT 148.630 10.500 155.490 13.500 ;
      LAYER li1 ;
        RECT 56.560 220.595 57.760 220.630 ;
        RECT 56.560 220.425 60.060 220.595 ;
        RECT 60.440 220.425 62.740 220.595 ;
        RECT 63.120 220.425 65.420 220.595 ;
        RECT 65.800 220.425 77.300 220.595 ;
        RECT 56.560 220.420 57.760 220.425 ;
        RECT 56.560 219.510 57.390 220.420 ;
        RECT 57.945 219.965 58.155 220.425 ;
        RECT 58.325 219.475 58.655 220.255 ;
        RECT 58.825 219.625 58.995 220.425 ;
        RECT 57.890 219.455 58.655 219.475 ;
        RECT 59.165 219.455 59.495 220.255 ;
        RECT 57.890 219.285 59.495 219.455 ;
        RECT 59.665 219.285 59.930 220.425 ;
        RECT 60.625 219.965 60.835 220.425 ;
        RECT 61.005 219.475 61.335 220.255 ;
        RECT 61.505 219.625 61.675 220.425 ;
        RECT 60.570 219.455 61.335 219.475 ;
        RECT 61.845 219.455 62.175 220.255 ;
        RECT 60.570 219.285 62.175 219.455 ;
        RECT 62.345 219.285 62.610 220.425 ;
        RECT 63.305 219.965 63.515 220.425 ;
        RECT 63.685 219.475 64.015 220.255 ;
        RECT 64.185 219.625 64.355 220.425 ;
        RECT 63.250 219.455 64.015 219.475 ;
        RECT 64.525 219.455 64.855 220.255 ;
        RECT 63.250 219.285 64.855 219.455 ;
        RECT 65.025 219.285 65.290 220.425 ;
        RECT 57.890 219.280 58.155 219.285 ;
        RECT 57.650 218.800 58.155 219.280 ;
        RECT 58.325 219.110 59.955 219.115 ;
        RECT 60.570 219.110 60.835 219.285 ;
        RECT 58.325 218.880 60.835 219.110 ;
        RECT 58.325 218.865 59.955 218.880 ;
        RECT 57.070 217.900 57.490 218.730 ;
        RECT 57.890 218.695 58.155 218.800 ;
        RECT 60.570 218.695 60.835 218.880 ;
        RECT 61.005 219.110 62.635 219.115 ;
        RECT 63.250 219.110 63.515 219.285 ;
        RECT 66.080 219.235 66.250 220.425 ;
        RECT 66.420 219.870 66.720 220.255 ;
        RECT 66.890 220.045 67.220 220.425 ;
        RECT 67.770 219.995 68.110 220.425 ;
        RECT 66.420 219.325 66.810 219.870 ;
        RECT 68.280 219.825 68.505 220.255 ;
        RECT 68.785 220.045 69.130 220.425 ;
        RECT 69.310 219.875 69.480 220.165 ;
        RECT 69.650 219.965 69.900 220.425 ;
        RECT 67.005 219.655 68.505 219.825 ;
        RECT 61.005 218.880 63.515 219.110 ;
        RECT 61.005 218.865 62.635 218.880 ;
        RECT 63.250 218.695 63.515 218.880 ;
        RECT 63.685 218.865 65.315 219.115 ;
        RECT 57.890 218.515 59.495 218.695 ;
        RECT 60.570 218.515 62.175 218.695 ;
        RECT 63.250 218.515 64.855 218.695 ;
        RECT 57.905 217.900 58.155 218.340 ;
        RECT 58.325 218.045 58.655 218.515 ;
        RECT 57.070 217.875 58.155 217.900 ;
        RECT 58.825 217.875 58.995 218.335 ;
        RECT 59.165 218.045 59.495 218.515 ;
        RECT 59.665 217.875 59.930 218.335 ;
        RECT 60.585 217.875 60.835 218.340 ;
        RECT 61.005 218.045 61.335 218.515 ;
        RECT 61.505 217.875 61.675 218.335 ;
        RECT 61.845 218.045 62.175 218.515 ;
        RECT 62.345 217.875 62.610 218.335 ;
        RECT 63.265 217.875 63.515 218.340 ;
        RECT 63.685 218.045 64.015 218.515 ;
        RECT 64.185 217.875 64.355 218.335 ;
        RECT 64.525 218.045 64.855 218.515 ;
        RECT 65.025 217.875 65.290 218.335 ;
        RECT 66.080 217.875 66.250 218.720 ;
        RECT 66.420 218.615 66.590 219.325 ;
        RECT 67.005 219.115 67.175 219.655 ;
        RECT 67.850 219.585 68.505 219.655 ;
        RECT 68.680 219.705 69.480 219.875 ;
        RECT 70.070 219.915 70.940 220.255 ;
        RECT 66.760 218.785 67.175 219.115 ;
        RECT 66.420 218.100 66.800 218.615 ;
        RECT 66.970 217.875 67.140 218.615 ;
        RECT 67.345 218.055 67.680 219.485 ;
        RECT 67.850 218.675 68.020 219.585 ;
        RECT 68.680 219.115 68.850 219.705 ;
        RECT 70.070 219.535 70.240 219.915 ;
        RECT 71.175 219.795 71.345 220.255 ;
        RECT 71.515 219.965 71.885 220.425 ;
        RECT 72.180 219.825 72.350 220.165 ;
        RECT 72.520 219.995 72.850 220.425 ;
        RECT 73.085 219.825 73.255 220.165 ;
        RECT 69.020 219.365 70.240 219.535 ;
        RECT 70.410 219.455 70.870 219.745 ;
        RECT 71.175 219.625 71.735 219.795 ;
        RECT 72.180 219.655 73.255 219.825 ;
        RECT 73.425 219.925 74.105 220.255 ;
        RECT 74.320 219.925 74.570 220.255 ;
        RECT 74.740 219.965 74.990 220.425 ;
        RECT 75.240 220.240 75.430 220.425 ;
        RECT 71.565 219.485 71.735 219.625 ;
        RECT 70.410 219.445 71.375 219.455 ;
        RECT 70.070 219.275 70.240 219.365 ;
        RECT 70.700 219.285 71.375 219.445 ;
        RECT 68.190 219.085 68.850 219.115 ;
        RECT 68.190 218.865 69.025 219.085 ;
        RECT 68.680 218.785 69.025 218.865 ;
        RECT 67.850 218.505 68.505 218.675 ;
        RECT 67.850 217.875 68.085 218.335 ;
        RECT 68.255 218.135 68.505 218.505 ;
        RECT 68.855 218.255 69.025 218.785 ;
        RECT 69.195 218.825 69.735 219.195 ;
        RECT 70.070 219.105 70.475 219.275 ;
        RECT 69.195 218.425 69.435 218.825 ;
        RECT 69.915 218.655 70.135 218.935 ;
        RECT 69.605 218.485 70.135 218.655 ;
        RECT 69.605 218.255 69.775 218.485 ;
        RECT 70.305 218.325 70.475 219.105 ;
        RECT 70.645 218.495 70.995 219.115 ;
        RECT 71.165 218.495 71.375 219.285 ;
        RECT 71.565 219.315 73.065 219.485 ;
        RECT 71.565 218.625 71.735 219.315 ;
        RECT 73.425 219.145 73.595 219.925 ;
        RECT 74.400 219.795 74.570 219.925 ;
        RECT 71.905 218.975 73.595 219.145 ;
        RECT 73.765 219.365 74.230 219.755 ;
        RECT 74.400 219.625 74.795 219.795 ;
        RECT 71.905 218.795 72.075 218.975 ;
        RECT 68.855 218.085 69.775 218.255 ;
        RECT 69.945 217.875 70.135 218.315 ;
        RECT 70.305 218.045 71.255 218.325 ;
        RECT 71.565 218.235 71.825 218.625 ;
        RECT 72.245 218.555 73.035 218.805 ;
        RECT 71.475 218.065 71.825 218.235 ;
        RECT 72.035 217.875 72.365 218.335 ;
        RECT 73.240 218.265 73.410 218.975 ;
        RECT 73.765 218.775 73.935 219.365 ;
        RECT 73.580 218.555 73.935 218.775 ;
        RECT 74.105 218.555 74.455 219.175 ;
        RECT 74.625 218.265 74.795 219.625 ;
        RECT 75.160 219.455 75.485 220.240 ;
        RECT 74.965 218.405 75.425 219.455 ;
        RECT 73.240 218.095 74.095 218.265 ;
        RECT 74.300 218.095 74.795 218.265 ;
        RECT 74.965 217.875 75.295 218.235 ;
        RECT 75.655 218.135 75.825 220.255 ;
        RECT 75.995 219.925 76.325 220.425 ;
        RECT 76.495 219.755 76.750 220.255 ;
        RECT 76.000 219.585 76.750 219.755 ;
        RECT 76.000 218.595 76.230 219.585 ;
        RECT 76.400 219.080 76.750 219.415 ;
        RECT 76.925 219.260 77.215 220.425 ;
        RECT 133.250 220.080 134.540 220.110 ;
        RECT 133.210 219.580 134.540 220.080 ;
        RECT 133.210 219.350 133.490 219.580 ;
        RECT 133.280 219.305 133.490 219.350 ;
        RECT 136.005 219.305 136.175 219.400 ;
        RECT 133.280 219.250 134.595 219.305 ;
        RECT 76.400 218.800 77.140 219.080 ;
        RECT 133.285 219.055 134.595 219.250 ;
        RECT 135.185 219.055 136.175 219.305 ;
        RECT 76.400 218.765 76.750 218.800 ;
        RECT 76.000 218.425 76.750 218.595 ;
        RECT 75.995 217.875 76.325 218.255 ;
        RECT 76.495 218.135 76.750 218.425 ;
        RECT 76.925 217.875 77.215 218.600 ;
        RECT 133.285 218.380 133.455 219.055 ;
        RECT 133.625 218.670 135.825 218.885 ;
        RECT 133.625 218.550 134.595 218.670 ;
        RECT 135.205 218.630 135.825 218.670 ;
        RECT 133.285 218.165 134.595 218.380 ;
        RECT 57.070 217.710 60.060 217.875 ;
        RECT 57.760 217.705 60.060 217.710 ;
        RECT 60.440 217.705 62.740 217.875 ;
        RECT 63.120 217.705 65.420 217.875 ;
        RECT 65.800 217.705 77.300 217.875 ;
        RECT 133.285 217.305 133.455 218.165 ;
        RECT 134.765 217.975 135.095 218.500 ;
        RECT 136.005 218.460 136.175 219.055 ;
        RECT 135.265 218.130 136.175 218.460 ;
        RECT 133.645 217.905 135.095 217.975 ;
        RECT 133.645 217.705 135.745 217.905 ;
        RECT 133.645 217.645 134.375 217.705 ;
        RECT 135.475 217.645 135.745 217.705 ;
        RECT 136.005 217.310 136.175 218.130 ;
        RECT 62.380 217.255 63.580 217.280 ;
        RECT 62.380 217.085 66.340 217.255 ;
        RECT 66.720 217.085 69.020 217.255 ;
        RECT 133.285 217.130 134.370 217.305 ;
        RECT 135.490 217.140 136.175 217.310 ;
        RECT 62.380 217.080 63.580 217.085 ;
        RECT 62.380 216.160 63.210 217.080 ;
        RECT 63.865 216.415 64.145 217.085 ;
        RECT 63.665 215.775 63.980 216.215 ;
        RECT 64.315 216.195 64.615 216.745 ;
        RECT 64.825 216.365 65.155 217.085 ;
        RECT 65.345 216.365 65.795 216.915 ;
        RECT 64.315 216.025 65.255 216.195 ;
        RECT 65.085 215.775 65.255 216.025 ;
        RECT 63.665 215.525 64.355 215.775 ;
        RECT 64.585 215.525 64.915 215.775 ;
        RECT 65.085 215.445 65.375 215.775 ;
        RECT 65.545 215.770 65.795 216.365 ;
        RECT 65.965 215.945 66.255 217.085 ;
        RECT 66.850 215.945 67.115 217.085 ;
        RECT 67.285 216.115 67.615 216.915 ;
        RECT 67.785 216.285 67.955 217.085 ;
        RECT 68.125 216.135 68.455 216.915 ;
        RECT 68.625 216.625 68.835 217.085 ;
        RECT 133.285 216.460 133.455 217.130 ;
        RECT 134.515 216.970 135.350 217.040 ;
        RECT 134.515 216.960 135.785 216.970 ;
        RECT 133.670 216.850 135.785 216.960 ;
        RECT 133.670 216.805 134.645 216.850 ;
        RECT 133.670 216.630 134.595 216.805 ;
        RECT 135.225 216.795 135.785 216.850 ;
        RECT 133.285 216.290 134.465 216.460 ;
        RECT 68.125 216.115 68.890 216.135 ;
        RECT 67.285 215.945 68.890 216.115 ;
        RECT 66.825 215.770 68.455 215.775 ;
        RECT 65.545 215.525 68.455 215.770 ;
        RECT 65.545 215.520 66.830 215.525 ;
        RECT 65.085 215.355 65.255 215.445 ;
        RECT 63.190 214.540 63.610 215.300 ;
        RECT 63.865 215.165 65.255 215.355 ;
        RECT 63.865 214.805 64.195 215.165 ;
        RECT 65.545 214.995 65.795 215.520 ;
        RECT 68.625 215.355 68.890 215.945 ;
        RECT 64.825 214.540 65.075 214.995 ;
        RECT 65.245 214.705 65.795 214.995 ;
        RECT 63.190 214.535 65.075 214.540 ;
        RECT 65.965 214.535 66.255 215.335 ;
        RECT 67.285 215.175 68.890 215.355 ;
        RECT 133.285 215.545 133.455 216.290 ;
        RECT 134.765 216.130 135.095 216.680 ;
        RECT 135.265 216.640 135.785 216.795 ;
        RECT 136.005 216.470 136.175 217.140 ;
        RECT 135.395 216.300 136.175 216.470 ;
        RECT 134.765 216.120 135.790 216.130 ;
        RECT 133.625 215.930 135.790 216.120 ;
        RECT 133.625 215.780 134.560 215.930 ;
        RECT 135.265 215.800 135.790 215.930 ;
        RECT 133.285 215.230 133.955 215.545 ;
        RECT 66.850 214.535 67.115 214.995 ;
        RECT 67.285 214.705 67.615 215.175 ;
        RECT 67.785 214.535 67.955 214.995 ;
        RECT 68.125 214.705 68.455 215.175 ;
        RECT 68.625 214.535 68.875 215.000 ;
        RECT 63.190 214.370 66.340 214.535 ;
        RECT 63.580 214.365 66.340 214.370 ;
        RECT 66.720 214.365 69.020 214.535 ;
        RECT 10.420 213.855 19.160 214.025 ;
        RECT 23.220 213.865 31.960 214.035 ;
        RECT 35.130 213.865 43.870 214.035 ;
        RECT 59.430 213.915 60.630 213.930 ;
        RECT 10.595 213.305 10.765 213.595 ;
        RECT 10.935 213.475 11.265 213.855 ;
        RECT 10.595 213.135 11.260 213.305 ;
        RECT 10.510 212.315 10.860 212.965 ;
        RECT 11.030 212.145 11.260 213.135 ;
        RECT 10.595 211.975 11.260 212.145 ;
        RECT 10.595 211.475 10.765 211.975 ;
        RECT 10.935 211.305 11.265 211.805 ;
        RECT 11.435 211.475 11.620 213.595 ;
        RECT 11.875 213.395 12.125 213.855 ;
        RECT 12.295 213.405 12.630 213.575 ;
        RECT 12.825 213.405 13.500 213.575 ;
        RECT 12.295 213.265 12.465 213.405 ;
        RECT 11.790 212.275 12.070 213.225 ;
        RECT 12.240 213.135 12.465 213.265 ;
        RECT 12.240 212.030 12.410 213.135 ;
        RECT 12.635 212.985 13.160 213.205 ;
        RECT 12.580 212.220 12.820 212.815 ;
        RECT 12.990 212.285 13.160 212.985 ;
        RECT 13.330 212.625 13.500 213.405 ;
        RECT 13.820 213.355 14.190 213.855 ;
        RECT 14.370 213.405 14.775 213.575 ;
        RECT 14.945 213.405 15.730 213.575 ;
        RECT 14.370 213.175 14.540 213.405 ;
        RECT 13.710 212.875 14.540 213.175 ;
        RECT 14.925 212.905 15.390 213.235 ;
        RECT 13.710 212.845 13.910 212.875 ;
        RECT 14.030 212.625 14.200 212.695 ;
        RECT 13.330 212.455 14.200 212.625 ;
        RECT 13.690 212.365 14.200 212.455 ;
        RECT 12.240 211.900 12.545 212.030 ;
        RECT 12.990 211.920 13.520 212.285 ;
        RECT 11.860 211.305 12.125 211.765 ;
        RECT 12.295 211.475 12.545 211.900 ;
        RECT 13.690 211.750 13.860 212.365 ;
        RECT 12.755 211.580 13.860 211.750 ;
        RECT 14.030 211.305 14.200 212.105 ;
        RECT 14.370 211.805 14.540 212.875 ;
        RECT 14.710 211.975 14.900 212.695 ;
        RECT 15.070 211.945 15.390 212.905 ;
        RECT 15.560 212.945 15.730 213.405 ;
        RECT 16.005 213.325 16.215 213.855 ;
        RECT 16.480 213.115 16.810 213.640 ;
        RECT 16.980 213.245 17.150 213.855 ;
        RECT 17.320 213.200 17.650 213.635 ;
        RECT 17.840 213.325 18.090 213.595 ;
        RECT 18.325 213.395 18.645 213.855 ;
        RECT 17.320 213.115 17.720 213.200 ;
        RECT 16.610 212.945 16.810 213.115 ;
        RECT 17.475 213.075 17.720 213.115 ;
        RECT 15.560 212.615 16.440 212.945 ;
        RECT 16.610 212.615 17.360 212.945 ;
        RECT 14.370 211.475 14.620 211.805 ;
        RECT 15.560 211.775 15.730 212.615 ;
        RECT 16.610 212.410 16.800 212.615 ;
        RECT 17.530 212.495 17.720 213.075 ;
        RECT 17.485 212.445 17.720 212.495 ;
        RECT 15.900 212.035 16.800 212.410 ;
        RECT 17.310 212.365 17.720 212.445 ;
        RECT 17.890 212.945 18.090 213.325 ;
        RECT 18.815 213.030 19.070 213.685 ;
        RECT 19.330 213.040 19.910 213.620 ;
        RECT 23.395 213.315 23.565 213.605 ;
        RECT 23.735 213.485 24.065 213.865 ;
        RECT 23.395 213.145 24.060 213.315 ;
        RECT 17.890 212.615 18.665 212.945 ;
        RECT 14.845 211.605 15.730 211.775 ;
        RECT 15.910 211.305 16.225 211.805 ;
        RECT 16.460 211.475 16.800 212.035 ;
        RECT 16.970 211.305 17.140 212.315 ;
        RECT 17.310 211.520 17.640 212.365 ;
        RECT 17.890 212.225 18.160 212.615 ;
        RECT 18.835 212.460 19.070 213.030 ;
        RECT 17.830 211.495 18.160 212.225 ;
        RECT 18.350 211.305 18.565 212.445 ;
        RECT 18.735 211.475 19.070 212.460 ;
        RECT 19.370 211.740 19.800 212.360 ;
        RECT 23.310 212.325 23.660 212.975 ;
        RECT 23.830 212.155 24.060 213.145 ;
        RECT 23.395 211.985 24.060 212.155 ;
        RECT 10.420 211.300 19.160 211.305 ;
        RECT 19.460 211.300 19.650 211.740 ;
        RECT 23.395 211.485 23.565 211.985 ;
        RECT 23.735 211.315 24.065 211.815 ;
        RECT 24.235 211.485 24.420 213.605 ;
        RECT 24.675 213.405 24.925 213.865 ;
        RECT 25.095 213.415 25.430 213.585 ;
        RECT 25.625 213.415 26.300 213.585 ;
        RECT 25.095 213.275 25.265 213.415 ;
        RECT 24.590 212.285 24.870 213.235 ;
        RECT 25.040 213.145 25.265 213.275 ;
        RECT 25.040 212.040 25.210 213.145 ;
        RECT 25.435 212.995 25.960 213.215 ;
        RECT 25.380 212.230 25.620 212.825 ;
        RECT 25.790 212.295 25.960 212.995 ;
        RECT 26.130 212.635 26.300 213.415 ;
        RECT 26.620 213.365 26.990 213.865 ;
        RECT 27.170 213.415 27.575 213.585 ;
        RECT 27.745 213.415 28.530 213.585 ;
        RECT 27.170 213.185 27.340 213.415 ;
        RECT 26.510 212.885 27.340 213.185 ;
        RECT 27.725 212.915 28.190 213.245 ;
        RECT 26.510 212.855 26.710 212.885 ;
        RECT 26.830 212.635 27.000 212.705 ;
        RECT 26.130 212.465 27.000 212.635 ;
        RECT 26.490 212.375 27.000 212.465 ;
        RECT 25.040 211.910 25.345 212.040 ;
        RECT 25.790 211.930 26.320 212.295 ;
        RECT 24.660 211.315 24.925 211.775 ;
        RECT 25.095 211.485 25.345 211.910 ;
        RECT 26.490 211.760 26.660 212.375 ;
        RECT 25.555 211.590 26.660 211.760 ;
        RECT 26.830 211.315 27.000 212.115 ;
        RECT 27.170 211.815 27.340 212.885 ;
        RECT 27.510 211.985 27.700 212.705 ;
        RECT 27.870 211.955 28.190 212.915 ;
        RECT 28.360 212.955 28.530 213.415 ;
        RECT 28.805 213.335 29.015 213.865 ;
        RECT 29.280 213.125 29.610 213.650 ;
        RECT 29.780 213.255 29.950 213.865 ;
        RECT 30.120 213.210 30.450 213.645 ;
        RECT 30.640 213.335 30.890 213.605 ;
        RECT 31.125 213.405 31.445 213.865 ;
        RECT 30.120 213.125 30.520 213.210 ;
        RECT 29.410 212.955 29.610 213.125 ;
        RECT 30.275 213.085 30.520 213.125 ;
        RECT 28.360 212.625 29.240 212.955 ;
        RECT 29.410 212.625 30.160 212.955 ;
        RECT 27.170 211.485 27.420 211.815 ;
        RECT 28.360 211.785 28.530 212.625 ;
        RECT 29.410 212.420 29.600 212.625 ;
        RECT 30.330 212.505 30.520 213.085 ;
        RECT 30.285 212.455 30.520 212.505 ;
        RECT 28.700 212.045 29.600 212.420 ;
        RECT 30.110 212.375 30.520 212.455 ;
        RECT 30.690 212.955 30.890 213.335 ;
        RECT 31.615 213.040 31.870 213.695 ;
        RECT 30.690 212.625 31.465 212.955 ;
        RECT 27.645 211.615 28.530 211.785 ;
        RECT 28.710 211.315 29.025 211.815 ;
        RECT 29.260 211.485 29.600 212.045 ;
        RECT 29.770 211.315 29.940 212.325 ;
        RECT 30.110 211.530 30.440 212.375 ;
        RECT 30.690 212.235 30.960 212.625 ;
        RECT 31.635 212.470 31.870 213.040 ;
        RECT 32.140 212.980 32.720 213.560 ;
        RECT 35.305 213.315 35.475 213.605 ;
        RECT 35.645 213.485 35.975 213.865 ;
        RECT 35.305 213.145 35.970 213.315 ;
        RECT 35.220 212.890 35.570 212.975 ;
        RECT 35.210 212.630 35.570 212.890 ;
        RECT 30.630 211.505 30.960 212.235 ;
        RECT 31.150 211.315 31.365 212.455 ;
        RECT 31.535 211.485 31.870 212.470 ;
        RECT 35.220 212.325 35.570 212.630 ;
        RECT 32.170 211.720 32.640 212.280 ;
        RECT 35.740 212.155 35.970 213.145 ;
        RECT 35.305 211.985 35.970 212.155 ;
        RECT 10.420 211.135 19.650 211.300 ;
        RECT 23.220 211.310 31.960 211.315 ;
        RECT 32.200 211.310 32.420 211.720 ;
        RECT 35.305 211.485 35.475 211.985 ;
        RECT 35.645 211.315 35.975 211.815 ;
        RECT 36.145 211.485 36.330 213.605 ;
        RECT 36.585 213.405 36.835 213.865 ;
        RECT 37.005 213.415 37.340 213.585 ;
        RECT 37.535 213.415 38.210 213.585 ;
        RECT 37.005 213.275 37.175 213.415 ;
        RECT 36.500 212.285 36.780 213.235 ;
        RECT 36.950 213.145 37.175 213.275 ;
        RECT 36.950 212.040 37.120 213.145 ;
        RECT 37.345 212.995 37.870 213.215 ;
        RECT 37.290 212.230 37.530 212.825 ;
        RECT 37.700 212.295 37.870 212.995 ;
        RECT 38.040 212.635 38.210 213.415 ;
        RECT 38.530 213.365 38.900 213.865 ;
        RECT 39.080 213.415 39.485 213.585 ;
        RECT 39.655 213.415 40.440 213.585 ;
        RECT 39.080 213.185 39.250 213.415 ;
        RECT 38.420 212.885 39.250 213.185 ;
        RECT 39.635 212.915 40.100 213.245 ;
        RECT 38.420 212.855 38.620 212.885 ;
        RECT 38.740 212.635 38.910 212.705 ;
        RECT 38.040 212.465 38.910 212.635 ;
        RECT 38.400 212.375 38.910 212.465 ;
        RECT 36.950 211.910 37.255 212.040 ;
        RECT 37.700 211.930 38.230 212.295 ;
        RECT 36.570 211.315 36.835 211.775 ;
        RECT 37.005 211.485 37.255 211.910 ;
        RECT 38.400 211.760 38.570 212.375 ;
        RECT 37.465 211.590 38.570 211.760 ;
        RECT 38.740 211.315 38.910 212.115 ;
        RECT 39.080 211.815 39.250 212.885 ;
        RECT 39.420 211.985 39.610 212.705 ;
        RECT 39.780 211.955 40.100 212.915 ;
        RECT 40.270 212.955 40.440 213.415 ;
        RECT 40.715 213.335 40.925 213.865 ;
        RECT 41.190 213.125 41.520 213.650 ;
        RECT 41.690 213.255 41.860 213.865 ;
        RECT 42.030 213.210 42.360 213.645 ;
        RECT 42.550 213.335 42.800 213.605 ;
        RECT 43.035 213.405 43.355 213.865 ;
        RECT 59.430 213.745 62.930 213.915 ;
        RECT 63.310 213.745 65.610 213.915 ;
        RECT 65.800 213.745 77.300 213.915 ;
        RECT 59.430 213.740 60.630 213.745 ;
        RECT 42.030 213.125 42.430 213.210 ;
        RECT 41.320 212.955 41.520 213.125 ;
        RECT 42.185 213.085 42.430 213.125 ;
        RECT 40.270 212.625 41.150 212.955 ;
        RECT 41.320 212.625 42.070 212.955 ;
        RECT 39.080 211.485 39.330 211.815 ;
        RECT 40.270 211.785 40.440 212.625 ;
        RECT 41.320 212.420 41.510 212.625 ;
        RECT 42.240 212.505 42.430 213.085 ;
        RECT 42.195 212.455 42.430 212.505 ;
        RECT 40.610 212.045 41.510 212.420 ;
        RECT 42.020 212.375 42.430 212.455 ;
        RECT 42.600 212.955 42.800 213.335 ;
        RECT 43.525 213.040 43.780 213.695 ;
        RECT 42.600 212.625 43.375 212.955 ;
        RECT 39.555 211.615 40.440 211.785 ;
        RECT 40.620 211.315 40.935 211.815 ;
        RECT 41.170 211.485 41.510 212.045 ;
        RECT 41.680 211.315 41.850 212.325 ;
        RECT 42.020 211.530 42.350 212.375 ;
        RECT 42.600 212.235 42.870 212.625 ;
        RECT 43.545 212.470 43.780 213.040 ;
        RECT 44.040 213.010 44.620 213.590 ;
        RECT 59.430 212.820 60.260 213.740 ;
        RECT 60.815 213.285 61.025 213.745 ;
        RECT 61.195 212.795 61.525 213.575 ;
        RECT 61.695 212.945 61.865 213.745 ;
        RECT 60.760 212.775 61.525 212.795 ;
        RECT 62.035 212.775 62.365 213.575 ;
        RECT 60.760 212.630 62.365 212.775 ;
        RECT 42.540 211.505 42.870 212.235 ;
        RECT 43.060 211.315 43.275 212.455 ;
        RECT 43.445 211.485 43.780 212.470 ;
        RECT 60.470 212.605 62.365 212.630 ;
        RECT 62.535 212.605 62.800 213.745 ;
        RECT 63.495 213.285 63.705 213.745 ;
        RECT 63.875 212.795 64.205 213.575 ;
        RECT 64.375 212.945 64.545 213.745 ;
        RECT 63.440 212.775 64.205 212.795 ;
        RECT 64.715 212.775 65.045 213.575 ;
        RECT 63.440 212.605 65.045 212.775 ;
        RECT 65.215 212.605 65.480 213.745 ;
        RECT 60.470 212.130 61.025 212.605 ;
        RECT 61.195 212.430 62.825 212.435 ;
        RECT 63.440 212.430 63.705 212.605 ;
        RECT 66.080 212.555 66.250 213.745 ;
        RECT 66.420 213.190 66.720 213.575 ;
        RECT 66.890 213.365 67.220 213.745 ;
        RECT 67.770 213.315 68.110 213.745 ;
        RECT 66.420 212.645 66.810 213.190 ;
        RECT 68.280 213.145 68.505 213.575 ;
        RECT 68.785 213.365 69.130 213.745 ;
        RECT 69.310 213.195 69.480 213.485 ;
        RECT 69.650 213.285 69.900 213.745 ;
        RECT 67.005 212.975 68.505 213.145 ;
        RECT 61.195 212.190 63.705 212.430 ;
        RECT 61.195 212.185 62.825 212.190 ;
        RECT 23.220 211.145 32.420 211.310 ;
        RECT 35.130 211.310 43.870 211.315 ;
        RECT 44.180 211.310 44.450 211.780 ;
        RECT 35.130 211.145 44.450 211.310 ;
        RECT 31.650 211.140 32.420 211.145 ;
        RECT 43.550 211.140 44.450 211.145 ;
        RECT 18.810 211.110 19.650 211.135 ;
        RECT 32.200 211.130 32.420 211.140 ;
        RECT 44.180 211.120 44.450 211.140 ;
        RECT 59.900 211.210 60.320 212.050 ;
        RECT 60.760 212.015 61.025 212.130 ;
        RECT 63.440 212.015 63.705 212.190 ;
        RECT 63.875 212.185 65.505 212.435 ;
        RECT 60.760 211.835 62.365 212.015 ;
        RECT 63.440 211.835 65.045 212.015 ;
        RECT 60.775 211.210 61.025 211.660 ;
        RECT 61.195 211.365 61.525 211.835 ;
        RECT 59.900 211.195 61.025 211.210 ;
        RECT 61.695 211.195 61.865 211.655 ;
        RECT 62.035 211.365 62.365 211.835 ;
        RECT 62.535 211.195 62.800 211.655 ;
        RECT 63.455 211.195 63.705 211.660 ;
        RECT 63.875 211.365 64.205 211.835 ;
        RECT 64.375 211.195 64.545 211.655 ;
        RECT 64.715 211.365 65.045 211.835 ;
        RECT 65.215 211.195 65.480 211.655 ;
        RECT 66.080 211.195 66.250 212.040 ;
        RECT 66.420 211.935 66.590 212.645 ;
        RECT 67.005 212.435 67.175 212.975 ;
        RECT 67.850 212.905 68.505 212.975 ;
        RECT 68.680 213.025 69.480 213.195 ;
        RECT 70.070 213.235 70.940 213.575 ;
        RECT 66.760 212.105 67.175 212.435 ;
        RECT 66.420 211.420 66.800 211.935 ;
        RECT 66.970 211.195 67.140 211.935 ;
        RECT 67.345 211.375 67.680 212.805 ;
        RECT 67.850 211.995 68.020 212.905 ;
        RECT 68.680 212.435 68.850 213.025 ;
        RECT 70.070 212.855 70.240 213.235 ;
        RECT 71.175 213.115 71.345 213.575 ;
        RECT 71.515 213.285 71.885 213.745 ;
        RECT 72.180 213.145 72.350 213.485 ;
        RECT 72.520 213.315 72.850 213.745 ;
        RECT 73.085 213.145 73.255 213.485 ;
        RECT 69.020 212.685 70.240 212.855 ;
        RECT 70.410 212.775 70.870 213.065 ;
        RECT 71.175 212.945 71.735 213.115 ;
        RECT 72.180 212.975 73.255 213.145 ;
        RECT 73.425 213.245 74.105 213.575 ;
        RECT 74.320 213.245 74.570 213.575 ;
        RECT 74.740 213.285 74.990 213.745 ;
        RECT 75.230 213.560 75.420 213.745 ;
        RECT 71.565 212.805 71.735 212.945 ;
        RECT 70.410 212.765 71.375 212.775 ;
        RECT 70.070 212.595 70.240 212.685 ;
        RECT 70.700 212.605 71.375 212.765 ;
        RECT 68.190 212.405 68.850 212.435 ;
        RECT 68.190 212.185 69.025 212.405 ;
        RECT 68.680 212.105 69.025 212.185 ;
        RECT 67.850 211.825 68.505 211.995 ;
        RECT 67.850 211.195 68.085 211.655 ;
        RECT 68.255 211.455 68.505 211.825 ;
        RECT 68.855 211.575 69.025 212.105 ;
        RECT 69.195 212.145 69.735 212.515 ;
        RECT 70.070 212.425 70.475 212.595 ;
        RECT 69.195 211.745 69.435 212.145 ;
        RECT 69.915 211.975 70.135 212.255 ;
        RECT 69.605 211.805 70.135 211.975 ;
        RECT 69.605 211.575 69.775 211.805 ;
        RECT 70.305 211.645 70.475 212.425 ;
        RECT 70.645 211.815 70.995 212.435 ;
        RECT 71.165 211.815 71.375 212.605 ;
        RECT 71.565 212.635 73.065 212.805 ;
        RECT 71.565 211.945 71.735 212.635 ;
        RECT 73.425 212.465 73.595 213.245 ;
        RECT 74.400 213.115 74.570 213.245 ;
        RECT 71.905 212.295 73.595 212.465 ;
        RECT 73.765 212.685 74.230 213.075 ;
        RECT 74.400 212.945 74.795 213.115 ;
        RECT 71.905 212.115 72.075 212.295 ;
        RECT 68.855 211.405 69.775 211.575 ;
        RECT 69.945 211.195 70.135 211.635 ;
        RECT 70.305 211.365 71.255 211.645 ;
        RECT 71.565 211.555 71.825 211.945 ;
        RECT 72.245 211.875 73.035 212.125 ;
        RECT 71.475 211.385 71.825 211.555 ;
        RECT 72.035 211.195 72.365 211.655 ;
        RECT 73.240 211.585 73.410 212.295 ;
        RECT 73.765 212.095 73.935 212.685 ;
        RECT 73.580 211.875 73.935 212.095 ;
        RECT 74.105 211.875 74.455 212.495 ;
        RECT 74.625 211.585 74.795 212.945 ;
        RECT 75.160 212.775 75.485 213.560 ;
        RECT 74.965 211.725 75.425 212.775 ;
        RECT 73.240 211.415 74.095 211.585 ;
        RECT 74.300 211.415 74.795 211.585 ;
        RECT 74.965 211.195 75.295 211.555 ;
        RECT 75.655 211.455 75.825 213.575 ;
        RECT 75.995 213.245 76.325 213.745 ;
        RECT 76.495 213.075 76.750 213.575 ;
        RECT 76.000 212.905 76.750 213.075 ;
        RECT 76.000 211.915 76.230 212.905 ;
        RECT 76.400 212.085 76.750 212.735 ;
        RECT 76.925 212.580 77.215 213.745 ;
        RECT 133.285 213.520 133.455 215.230 ;
        RECT 134.185 215.220 134.560 215.780 ;
        RECT 134.765 215.050 135.095 215.760 ;
        RECT 136.005 215.535 136.175 216.300 ;
        RECT 135.475 215.325 136.175 215.535 ;
        RECT 133.755 214.880 135.725 215.050 ;
        RECT 133.755 214.165 133.925 214.880 ;
        RECT 134.095 214.390 135.385 214.710 ;
        RECT 135.055 214.245 135.385 214.390 ;
        RECT 135.555 214.265 135.725 214.880 ;
        RECT 134.125 214.030 134.845 214.220 ;
        RECT 133.625 213.860 133.955 213.940 ;
        RECT 135.555 213.860 135.725 214.095 ;
        RECT 133.625 213.690 135.725 213.860 ;
        RECT 133.285 213.350 134.255 213.520 ;
        RECT 134.515 213.350 134.845 213.520 ;
        RECT 76.000 211.745 76.750 211.915 ;
        RECT 75.995 211.195 76.325 211.575 ;
        RECT 76.495 211.455 76.750 211.745 ;
        RECT 76.925 211.195 77.215 211.920 ;
        RECT 133.285 211.445 133.455 213.350 ;
        RECT 134.515 213.180 134.775 213.350 ;
        RECT 135.025 213.230 135.325 213.690 ;
        RECT 136.005 213.510 136.175 215.325 ;
        RECT 133.730 213.010 134.775 213.180 ;
        RECT 134.995 213.030 135.325 213.230 ;
        RECT 135.505 213.140 136.175 213.510 ;
        RECT 133.730 212.075 133.900 213.010 ;
        RECT 134.070 212.480 134.435 212.840 ;
        RECT 134.605 212.820 134.775 213.010 ;
        RECT 134.605 212.650 135.725 212.820 ;
        RECT 134.070 212.310 135.355 212.480 ;
        RECT 134.370 211.900 134.965 212.140 ;
        RECT 135.135 211.955 135.355 212.310 ;
        RECT 135.555 212.145 135.725 212.650 ;
        RECT 133.625 211.730 134.180 211.865 ;
        RECT 135.555 211.785 135.725 211.950 ;
        RECT 135.285 211.730 135.725 211.785 ;
        RECT 133.625 211.615 135.725 211.730 ;
        RECT 134.050 211.560 135.415 211.615 ;
        RECT 136.005 211.445 136.175 213.140 ;
        RECT 59.900 211.030 62.930 211.195 ;
        RECT 60.630 211.025 62.930 211.030 ;
        RECT 63.310 211.025 65.610 211.195 ;
        RECT 65.800 211.025 77.300 211.195 ;
        RECT 133.285 211.180 133.915 211.445 ;
        RECT 133.285 210.585 133.455 211.180 ;
        RECT 134.425 211.110 135.375 211.390 ;
        RECT 135.545 211.195 136.175 211.445 ;
        RECT 133.625 210.755 135.745 210.940 ;
        RECT 136.005 210.585 136.175 211.195 ;
        RECT 133.285 210.255 133.955 210.585 ;
        RECT 134.125 210.350 135.455 210.580 ;
        RECT 133.285 209.655 133.455 210.255 ;
        RECT 134.125 210.085 134.295 210.350 ;
        RECT 133.625 209.915 134.295 210.085 ;
        RECT 134.465 209.830 135.115 210.180 ;
        RECT 135.285 210.085 135.455 210.350 ;
        RECT 135.625 210.255 136.175 210.585 ;
        RECT 135.285 209.915 135.745 210.085 ;
        RECT 133.285 209.365 134.620 209.655 ;
        RECT 133.285 209.185 133.455 209.365 ;
        RECT 133.285 208.935 134.595 209.185 ;
        RECT 133.285 208.260 133.455 208.935 ;
        RECT 134.820 208.765 134.990 209.830 ;
        RECT 136.005 209.655 136.175 210.255 ;
        RECT 135.280 209.365 136.175 209.655 ;
        RECT 136.005 209.185 136.175 209.365 ;
        RECT 135.185 208.935 136.175 209.185 ;
        RECT 133.625 208.550 135.825 208.765 ;
        RECT 133.625 208.430 134.595 208.550 ;
        RECT 135.205 208.510 135.825 208.550 ;
        RECT 133.285 208.045 134.595 208.260 ;
        RECT 133.285 207.185 133.455 208.045 ;
        RECT 134.765 207.855 135.095 208.380 ;
        RECT 136.005 208.340 136.175 208.935 ;
        RECT 135.265 208.010 136.175 208.340 ;
        RECT 133.645 207.785 135.095 207.855 ;
        RECT 133.645 207.585 135.745 207.785 ;
        RECT 133.645 207.525 134.375 207.585 ;
        RECT 135.475 207.525 135.745 207.585 ;
        RECT 136.005 207.190 136.175 208.010 ;
        RECT 133.285 207.010 134.370 207.185 ;
        RECT 135.490 207.020 136.175 207.190 ;
        RECT 133.285 206.340 133.455 207.010 ;
        RECT 134.515 206.850 135.350 206.920 ;
        RECT 134.515 206.840 135.785 206.850 ;
        RECT 133.670 206.730 135.785 206.840 ;
        RECT 133.670 206.685 134.645 206.730 ;
        RECT 133.670 206.510 134.595 206.685 ;
        RECT 135.225 206.675 135.785 206.730 ;
        RECT 85.640 206.020 86.150 206.180 ;
        RECT 133.285 206.170 134.465 206.340 ;
        RECT 85.640 205.830 87.970 206.020 ;
        RECT 85.640 205.140 86.150 205.830 ;
        RECT 86.590 205.825 87.970 205.830 ;
        RECT 88.160 205.825 89.540 205.995 ;
        RECT 89.770 205.825 98.510 205.995 ;
        RECT 98.700 205.825 99.160 205.995 ;
        RECT 99.370 205.825 108.110 205.995 ;
        RECT 108.280 205.825 117.480 205.995 ;
        RECT 86.735 204.685 86.945 205.825 ;
        RECT 87.115 204.675 87.445 205.655 ;
        RECT 87.615 204.685 87.845 205.825 ;
        RECT 88.305 204.685 88.515 205.825 ;
        RECT 88.685 204.675 89.015 205.655 ;
        RECT 89.185 204.685 89.415 205.825 ;
        RECT 86.320 204.500 86.570 204.620 ;
        RECT 87.115 204.500 87.365 204.675 ;
        RECT 86.320 204.300 87.365 204.500 ;
        RECT 86.320 204.170 86.570 204.300 ;
        RECT 85.650 203.340 86.140 204.130 ;
        RECT 86.735 203.340 86.945 204.095 ;
        RECT 87.115 204.075 87.365 204.300 ;
        RECT 87.535 204.510 87.865 204.515 ;
        RECT 88.685 204.510 88.935 204.675 ;
        RECT 89.860 204.670 90.195 205.655 ;
        RECT 90.365 204.685 90.580 205.825 ;
        RECT 90.770 204.905 91.100 205.635 ;
        RECT 87.535 204.270 88.935 204.510 ;
        RECT 87.535 204.265 87.865 204.270 ;
        RECT 87.115 203.445 87.445 204.075 ;
        RECT 85.650 203.275 86.945 203.340 ;
        RECT 87.615 203.275 87.845 204.095 ;
        RECT 88.305 203.275 88.515 204.095 ;
        RECT 88.685 204.075 88.935 204.270 ;
        RECT 89.105 204.265 89.435 204.515 ;
        RECT 89.860 204.100 90.095 204.670 ;
        RECT 90.770 204.515 91.040 204.905 ;
        RECT 91.290 204.765 91.620 205.610 ;
        RECT 91.790 204.815 91.960 205.825 ;
        RECT 92.130 205.095 92.470 205.655 ;
        RECT 92.705 205.325 93.020 205.825 ;
        RECT 93.200 205.355 94.085 205.525 ;
        RECT 90.265 204.185 91.040 204.515 ;
        RECT 88.685 203.445 89.015 204.075 ;
        RECT 89.185 203.275 89.415 204.095 ;
        RECT 89.860 203.445 90.115 204.100 ;
        RECT 90.840 203.805 91.040 204.185 ;
        RECT 91.210 204.685 91.620 204.765 ;
        RECT 92.130 204.720 93.030 205.095 ;
        RECT 91.210 204.635 91.445 204.685 ;
        RECT 91.210 204.055 91.400 204.635 ;
        RECT 92.130 204.515 92.320 204.720 ;
        RECT 93.200 204.515 93.370 205.355 ;
        RECT 94.310 205.325 94.560 205.655 ;
        RECT 91.570 204.185 92.320 204.515 ;
        RECT 92.490 204.185 93.370 204.515 ;
        RECT 91.210 204.015 91.455 204.055 ;
        RECT 92.120 204.015 92.320 204.185 ;
        RECT 91.210 203.930 91.610 204.015 ;
        RECT 90.285 203.275 90.605 203.735 ;
        RECT 90.840 203.535 91.090 203.805 ;
        RECT 91.280 203.495 91.610 203.930 ;
        RECT 91.780 203.275 91.950 203.885 ;
        RECT 92.120 203.490 92.450 204.015 ;
        RECT 92.715 203.275 92.925 203.805 ;
        RECT 93.200 203.725 93.370 204.185 ;
        RECT 93.540 204.225 93.860 205.185 ;
        RECT 94.030 204.435 94.220 205.155 ;
        RECT 94.390 204.255 94.560 205.325 ;
        RECT 94.730 205.025 94.900 205.825 ;
        RECT 95.070 205.380 96.175 205.550 ;
        RECT 95.070 204.765 95.240 205.380 ;
        RECT 96.385 205.230 96.635 205.655 ;
        RECT 96.805 205.365 97.070 205.825 ;
        RECT 95.410 204.845 95.940 205.210 ;
        RECT 96.385 205.100 96.690 205.230 ;
        RECT 94.730 204.675 95.240 204.765 ;
        RECT 94.730 204.505 95.600 204.675 ;
        RECT 94.730 204.435 94.900 204.505 ;
        RECT 95.020 204.255 95.220 204.285 ;
        RECT 93.540 203.895 94.005 204.225 ;
        RECT 94.390 203.955 95.220 204.255 ;
        RECT 94.390 203.725 94.560 203.955 ;
        RECT 93.200 203.555 93.985 203.725 ;
        RECT 94.155 203.555 94.560 203.725 ;
        RECT 94.740 203.275 95.110 203.775 ;
        RECT 95.430 203.725 95.600 204.505 ;
        RECT 95.770 204.145 95.940 204.845 ;
        RECT 96.110 204.315 96.350 204.910 ;
        RECT 95.770 203.925 96.295 204.145 ;
        RECT 96.520 203.995 96.690 205.100 ;
        RECT 96.465 203.865 96.690 203.995 ;
        RECT 96.860 203.905 97.140 204.855 ;
        RECT 96.465 203.725 96.635 203.865 ;
        RECT 95.430 203.555 96.105 203.725 ;
        RECT 96.300 203.555 96.635 203.725 ;
        RECT 96.805 203.275 97.055 203.735 ;
        RECT 97.310 203.535 97.495 205.655 ;
        RECT 97.665 205.325 97.995 205.825 ;
        RECT 98.165 205.155 98.335 205.655 ;
        RECT 97.670 204.985 98.335 205.155 ;
        RECT 97.670 203.995 97.900 204.985 ;
        RECT 98.070 204.480 98.420 204.815 ;
        RECT 98.785 204.660 99.075 205.825 ;
        RECT 99.460 204.670 99.795 205.655 ;
        RECT 99.965 204.685 100.180 205.825 ;
        RECT 100.370 204.905 100.700 205.635 ;
        RECT 99.460 204.480 99.695 204.670 ;
        RECT 100.370 204.515 100.640 204.905 ;
        RECT 100.890 204.765 101.220 205.610 ;
        RECT 101.390 204.815 101.560 205.825 ;
        RECT 101.730 205.095 102.070 205.655 ;
        RECT 102.305 205.325 102.620 205.825 ;
        RECT 102.800 205.355 103.685 205.525 ;
        RECT 98.070 204.200 99.695 204.480 ;
        RECT 98.070 204.165 98.420 204.200 ;
        RECT 99.460 204.100 99.695 204.200 ;
        RECT 99.865 204.185 100.640 204.515 ;
        RECT 97.670 203.825 98.335 203.995 ;
        RECT 97.665 203.275 97.995 203.655 ;
        RECT 98.165 203.535 98.335 203.825 ;
        RECT 98.785 203.275 99.075 204.000 ;
        RECT 99.460 203.445 99.715 204.100 ;
        RECT 100.440 203.805 100.640 204.185 ;
        RECT 100.810 204.685 101.220 204.765 ;
        RECT 101.730 204.720 102.630 205.095 ;
        RECT 100.810 204.635 101.045 204.685 ;
        RECT 100.810 204.055 101.000 204.635 ;
        RECT 101.730 204.515 101.920 204.720 ;
        RECT 102.800 204.515 102.970 205.355 ;
        RECT 103.910 205.325 104.160 205.655 ;
        RECT 101.170 204.185 101.920 204.515 ;
        RECT 102.090 204.185 102.970 204.515 ;
        RECT 100.810 204.015 101.055 204.055 ;
        RECT 101.720 204.015 101.920 204.185 ;
        RECT 100.810 203.930 101.210 204.015 ;
        RECT 99.885 203.275 100.205 203.735 ;
        RECT 100.440 203.535 100.690 203.805 ;
        RECT 100.880 203.495 101.210 203.930 ;
        RECT 101.380 203.275 101.550 203.885 ;
        RECT 101.720 203.490 102.050 204.015 ;
        RECT 102.315 203.275 102.525 203.805 ;
        RECT 102.800 203.725 102.970 204.185 ;
        RECT 103.140 204.225 103.460 205.185 ;
        RECT 103.630 204.435 103.820 205.155 ;
        RECT 103.990 204.255 104.160 205.325 ;
        RECT 104.330 205.025 104.500 205.825 ;
        RECT 104.670 205.380 105.775 205.550 ;
        RECT 104.670 204.765 104.840 205.380 ;
        RECT 105.985 205.230 106.235 205.655 ;
        RECT 106.405 205.365 106.670 205.825 ;
        RECT 105.010 204.845 105.540 205.210 ;
        RECT 105.985 205.100 106.290 205.230 ;
        RECT 104.330 204.675 104.840 204.765 ;
        RECT 104.330 204.505 105.200 204.675 ;
        RECT 104.330 204.435 104.500 204.505 ;
        RECT 104.620 204.255 104.820 204.285 ;
        RECT 103.140 203.895 103.605 204.225 ;
        RECT 103.990 203.955 104.820 204.255 ;
        RECT 103.990 203.725 104.160 203.955 ;
        RECT 102.800 203.555 103.585 203.725 ;
        RECT 103.755 203.555 104.160 203.725 ;
        RECT 104.340 203.275 104.710 203.775 ;
        RECT 105.030 203.725 105.200 204.505 ;
        RECT 105.370 204.145 105.540 204.845 ;
        RECT 105.710 204.315 105.950 204.910 ;
        RECT 105.370 203.925 105.895 204.145 ;
        RECT 106.120 203.995 106.290 205.100 ;
        RECT 106.065 203.865 106.290 203.995 ;
        RECT 106.460 203.905 106.740 204.855 ;
        RECT 106.065 203.725 106.235 203.865 ;
        RECT 105.030 203.555 105.705 203.725 ;
        RECT 105.900 203.555 106.235 203.725 ;
        RECT 106.405 203.275 106.655 203.735 ;
        RECT 106.910 203.535 107.095 205.655 ;
        RECT 107.265 205.325 107.595 205.825 ;
        RECT 107.765 205.155 107.935 205.655 ;
        RECT 107.270 204.985 107.935 205.155 ;
        RECT 107.270 203.995 107.500 204.985 ;
        RECT 107.670 204.790 108.020 204.815 ;
        RECT 108.370 204.790 108.705 205.655 ;
        RECT 107.670 204.670 108.705 204.790 ;
        RECT 108.875 204.685 109.090 205.825 ;
        RECT 109.280 204.905 109.610 205.635 ;
        RECT 107.670 204.460 108.605 204.670 ;
        RECT 109.280 204.515 109.550 204.905 ;
        RECT 109.800 204.765 110.130 205.610 ;
        RECT 110.300 204.815 110.470 205.825 ;
        RECT 110.640 205.095 110.980 205.655 ;
        RECT 111.215 205.325 111.530 205.825 ;
        RECT 111.710 205.355 112.595 205.525 ;
        RECT 107.670 204.165 108.020 204.460 ;
        RECT 108.370 204.100 108.605 204.460 ;
        RECT 108.775 204.185 109.550 204.515 ;
        RECT 107.270 203.825 107.935 203.995 ;
        RECT 107.265 203.275 107.595 203.655 ;
        RECT 107.765 203.535 107.935 203.825 ;
        RECT 108.370 203.445 108.625 204.100 ;
        RECT 109.350 203.805 109.550 204.185 ;
        RECT 109.720 204.685 110.130 204.765 ;
        RECT 110.640 204.720 111.540 205.095 ;
        RECT 109.720 204.635 109.955 204.685 ;
        RECT 109.720 204.055 109.910 204.635 ;
        RECT 110.640 204.515 110.830 204.720 ;
        RECT 111.710 204.515 111.880 205.355 ;
        RECT 112.820 205.325 113.070 205.655 ;
        RECT 110.080 204.185 110.830 204.515 ;
        RECT 111.000 204.185 111.880 204.515 ;
        RECT 109.720 204.015 109.965 204.055 ;
        RECT 110.630 204.015 110.830 204.185 ;
        RECT 109.720 203.930 110.120 204.015 ;
        RECT 108.795 203.275 109.115 203.735 ;
        RECT 109.350 203.535 109.600 203.805 ;
        RECT 109.790 203.495 110.120 203.930 ;
        RECT 110.290 203.275 110.460 203.885 ;
        RECT 110.630 203.490 110.960 204.015 ;
        RECT 111.225 203.275 111.435 203.805 ;
        RECT 111.710 203.725 111.880 204.185 ;
        RECT 112.050 204.225 112.370 205.185 ;
        RECT 112.540 204.435 112.730 205.155 ;
        RECT 112.900 204.255 113.070 205.325 ;
        RECT 113.240 205.025 113.410 205.825 ;
        RECT 113.580 205.380 114.685 205.550 ;
        RECT 113.580 204.765 113.750 205.380 ;
        RECT 114.895 205.230 115.145 205.655 ;
        RECT 115.315 205.365 115.580 205.825 ;
        RECT 113.920 204.845 114.450 205.210 ;
        RECT 114.895 205.100 115.200 205.230 ;
        RECT 113.240 204.675 113.750 204.765 ;
        RECT 113.240 204.505 114.110 204.675 ;
        RECT 113.240 204.435 113.410 204.505 ;
        RECT 113.530 204.255 113.730 204.285 ;
        RECT 112.050 203.895 112.515 204.225 ;
        RECT 112.900 203.955 113.730 204.255 ;
        RECT 112.900 203.725 113.070 203.955 ;
        RECT 111.710 203.555 112.495 203.725 ;
        RECT 112.665 203.555 113.070 203.725 ;
        RECT 113.250 203.275 113.620 203.775 ;
        RECT 113.940 203.725 114.110 204.505 ;
        RECT 114.280 204.145 114.450 204.845 ;
        RECT 114.620 204.315 114.860 204.910 ;
        RECT 114.280 203.925 114.805 204.145 ;
        RECT 115.030 203.995 115.200 205.100 ;
        RECT 114.975 203.865 115.200 203.995 ;
        RECT 115.370 203.905 115.650 204.855 ;
        RECT 114.975 203.725 115.145 203.865 ;
        RECT 113.940 203.555 114.615 203.725 ;
        RECT 114.810 203.555 115.145 203.725 ;
        RECT 115.315 203.275 115.565 203.735 ;
        RECT 115.820 203.535 116.005 205.655 ;
        RECT 116.175 205.325 116.505 205.825 ;
        RECT 116.675 205.155 116.845 205.655 ;
        RECT 116.180 204.985 116.845 205.155 ;
        RECT 116.180 203.995 116.410 204.985 ;
        RECT 116.580 204.360 116.930 204.815 ;
        RECT 117.105 204.660 117.395 205.825 ;
        RECT 133.285 205.425 133.455 206.170 ;
        RECT 134.765 206.010 135.095 206.560 ;
        RECT 135.265 206.520 135.785 206.675 ;
        RECT 136.005 206.350 136.175 207.020 ;
        RECT 135.395 206.180 136.175 206.350 ;
        RECT 134.765 206.000 135.790 206.010 ;
        RECT 133.625 205.810 135.790 206.000 ;
        RECT 133.625 205.660 134.560 205.810 ;
        RECT 135.265 205.680 135.790 205.810 ;
        RECT 133.285 205.110 133.955 205.425 ;
        RECT 116.580 204.190 117.510 204.360 ;
        RECT 116.580 204.165 116.930 204.190 ;
        RECT 116.180 203.825 116.845 203.995 ;
        RECT 116.175 203.275 116.505 203.655 ;
        RECT 116.675 203.535 116.845 203.825 ;
        RECT 117.105 203.275 117.395 204.000 ;
        RECT 133.285 203.400 133.455 205.110 ;
        RECT 134.185 205.100 134.560 205.660 ;
        RECT 134.765 204.930 135.095 205.640 ;
        RECT 136.005 205.415 136.175 206.180 ;
        RECT 135.475 205.205 136.175 205.415 ;
        RECT 133.755 204.760 135.725 204.930 ;
        RECT 133.755 204.045 133.925 204.760 ;
        RECT 134.095 204.270 135.385 204.590 ;
        RECT 135.055 204.125 135.385 204.270 ;
        RECT 135.555 204.145 135.725 204.760 ;
        RECT 134.125 203.910 134.845 204.100 ;
        RECT 133.625 203.740 133.955 203.820 ;
        RECT 135.555 203.740 135.725 203.975 ;
        RECT 133.625 203.570 135.725 203.740 ;
        RECT 85.650 203.110 87.970 203.275 ;
        RECT 86.590 203.105 87.970 203.110 ;
        RECT 88.160 203.105 89.540 203.275 ;
        RECT 89.770 203.105 98.510 203.275 ;
        RECT 98.700 203.105 99.160 203.275 ;
        RECT 99.370 203.105 108.110 203.275 ;
        RECT 108.280 203.105 117.480 203.275 ;
        RECT 133.285 203.230 134.255 203.400 ;
        RECT 134.515 203.230 134.845 203.400 ;
        RECT 20.480 202.465 20.800 202.470 ;
        RECT 11.140 202.295 20.800 202.465 ;
        RECT 23.560 202.295 33.220 202.465 ;
        RECT 11.315 201.625 11.485 202.125 ;
        RECT 11.655 201.795 11.985 202.295 ;
        RECT 11.315 201.455 11.980 201.625 ;
        RECT 11.230 200.635 11.580 201.285 ;
        RECT 11.750 200.465 11.980 201.455 ;
        RECT 11.315 200.295 11.980 200.465 ;
        RECT 11.315 200.005 11.485 200.295 ;
        RECT 11.655 199.745 11.985 200.125 ;
        RECT 12.155 200.005 12.340 202.125 ;
        RECT 12.580 201.835 12.845 202.295 ;
        RECT 13.015 201.700 13.265 202.125 ;
        RECT 13.475 201.850 14.580 202.020 ;
        RECT 12.960 201.570 13.265 201.700 ;
        RECT 12.510 200.375 12.790 201.325 ;
        RECT 12.960 200.465 13.130 201.570 ;
        RECT 13.300 200.785 13.540 201.380 ;
        RECT 13.710 201.315 14.240 201.680 ;
        RECT 13.710 200.615 13.880 201.315 ;
        RECT 14.410 201.235 14.580 201.850 ;
        RECT 14.750 201.495 14.920 202.295 ;
        RECT 15.090 201.795 15.340 202.125 ;
        RECT 15.565 201.825 16.450 201.995 ;
        RECT 14.410 201.145 14.920 201.235 ;
        RECT 12.960 200.335 13.185 200.465 ;
        RECT 13.355 200.395 13.880 200.615 ;
        RECT 14.050 200.975 14.920 201.145 ;
        RECT 12.595 199.745 12.845 200.205 ;
        RECT 13.015 200.195 13.185 200.335 ;
        RECT 14.050 200.195 14.220 200.975 ;
        RECT 14.750 200.905 14.920 200.975 ;
        RECT 14.430 200.725 14.630 200.755 ;
        RECT 15.090 200.725 15.260 201.795 ;
        RECT 15.430 200.905 15.620 201.625 ;
        RECT 14.430 200.425 15.260 200.725 ;
        RECT 15.790 200.695 16.110 201.655 ;
        RECT 13.015 200.025 13.350 200.195 ;
        RECT 13.545 200.025 14.220 200.195 ;
        RECT 14.540 199.745 14.910 200.245 ;
        RECT 15.090 200.195 15.260 200.425 ;
        RECT 15.645 200.365 16.110 200.695 ;
        RECT 16.280 200.985 16.450 201.825 ;
        RECT 16.630 201.795 16.945 202.295 ;
        RECT 17.180 201.565 17.520 202.125 ;
        RECT 16.620 201.190 17.520 201.565 ;
        RECT 17.690 201.285 17.860 202.295 ;
        RECT 17.330 200.985 17.520 201.190 ;
        RECT 18.030 201.235 18.360 202.080 ;
        RECT 18.530 201.380 18.705 202.295 ;
        RECT 19.045 201.375 19.375 202.105 ;
        RECT 18.030 201.155 18.440 201.235 ;
        RECT 18.205 201.105 18.440 201.155 ;
        RECT 16.280 200.655 17.160 200.985 ;
        RECT 17.330 200.655 18.080 200.985 ;
        RECT 16.280 200.195 16.450 200.655 ;
        RECT 17.330 200.485 17.530 200.655 ;
        RECT 18.250 200.525 18.440 201.105 ;
        RECT 18.195 200.485 18.440 200.525 ;
        RECT 15.090 200.025 15.495 200.195 ;
        RECT 15.665 200.025 16.450 200.195 ;
        RECT 16.725 199.745 16.935 200.275 ;
        RECT 17.200 199.960 17.530 200.485 ;
        RECT 18.040 200.400 18.440 200.485 ;
        RECT 19.105 200.985 19.375 201.375 ;
        RECT 19.565 201.155 19.780 202.295 ;
        RECT 20.455 202.260 20.800 202.295 ;
        RECT 19.950 201.155 20.285 202.125 ;
        RECT 20.455 202.000 21.360 202.260 ;
        RECT 20.455 201.155 20.705 202.000 ;
        RECT 23.735 201.625 23.905 202.125 ;
        RECT 24.075 201.795 24.405 202.295 ;
        RECT 23.735 201.455 24.400 201.625 ;
        RECT 19.105 200.655 19.900 200.985 ;
        RECT 17.700 199.745 17.870 200.355 ;
        RECT 18.040 199.965 18.370 200.400 ;
        RECT 19.105 200.275 19.305 200.655 ;
        RECT 20.070 200.545 20.285 201.155 ;
        RECT 23.650 200.635 24.000 201.285 ;
        RECT 18.540 199.745 18.710 200.260 ;
        RECT 19.045 200.005 19.305 200.275 ;
        RECT 19.530 199.745 19.860 200.485 ;
        RECT 20.030 199.925 20.285 200.545 ;
        RECT 20.455 200.470 20.705 200.565 ;
        RECT 20.455 200.230 21.410 200.470 ;
        RECT 24.170 200.465 24.400 201.455 ;
        RECT 23.735 200.295 24.400 200.465 ;
        RECT 20.455 199.745 20.705 200.230 ;
        RECT 23.735 200.005 23.905 200.295 ;
        RECT 24.075 199.745 24.405 200.125 ;
        RECT 24.575 200.005 24.760 202.125 ;
        RECT 25.000 201.835 25.265 202.295 ;
        RECT 25.435 201.700 25.685 202.125 ;
        RECT 25.895 201.850 27.000 202.020 ;
        RECT 25.380 201.570 25.685 201.700 ;
        RECT 24.930 200.375 25.210 201.325 ;
        RECT 25.380 200.465 25.550 201.570 ;
        RECT 25.720 200.785 25.960 201.380 ;
        RECT 26.130 201.315 26.660 201.680 ;
        RECT 26.130 200.615 26.300 201.315 ;
        RECT 26.830 201.235 27.000 201.850 ;
        RECT 27.170 201.495 27.340 202.295 ;
        RECT 27.510 201.795 27.760 202.125 ;
        RECT 27.985 201.825 28.870 201.995 ;
        RECT 26.830 201.145 27.340 201.235 ;
        RECT 25.380 200.335 25.605 200.465 ;
        RECT 25.775 200.395 26.300 200.615 ;
        RECT 26.470 200.975 27.340 201.145 ;
        RECT 25.015 199.745 25.265 200.205 ;
        RECT 25.435 200.195 25.605 200.335 ;
        RECT 26.470 200.195 26.640 200.975 ;
        RECT 27.170 200.905 27.340 200.975 ;
        RECT 26.850 200.725 27.050 200.755 ;
        RECT 27.510 200.725 27.680 201.795 ;
        RECT 27.850 200.905 28.040 201.625 ;
        RECT 26.850 200.425 27.680 200.725 ;
        RECT 28.210 200.695 28.530 201.655 ;
        RECT 25.435 200.025 25.770 200.195 ;
        RECT 25.965 200.025 26.640 200.195 ;
        RECT 26.960 199.745 27.330 200.245 ;
        RECT 27.510 200.195 27.680 200.425 ;
        RECT 28.065 200.365 28.530 200.695 ;
        RECT 28.700 200.985 28.870 201.825 ;
        RECT 29.050 201.795 29.365 202.295 ;
        RECT 29.600 201.565 29.940 202.125 ;
        RECT 29.040 201.190 29.940 201.565 ;
        RECT 30.110 201.285 30.280 202.295 ;
        RECT 29.750 200.985 29.940 201.190 ;
        RECT 30.450 201.235 30.780 202.080 ;
        RECT 30.950 201.380 31.125 202.295 ;
        RECT 31.465 201.375 31.795 202.105 ;
        RECT 30.450 201.155 30.860 201.235 ;
        RECT 30.625 201.105 30.860 201.155 ;
        RECT 28.700 200.655 29.580 200.985 ;
        RECT 29.750 200.655 30.500 200.985 ;
        RECT 28.700 200.195 28.870 200.655 ;
        RECT 29.750 200.485 29.950 200.655 ;
        RECT 30.670 200.525 30.860 201.105 ;
        RECT 30.615 200.485 30.860 200.525 ;
        RECT 27.510 200.025 27.915 200.195 ;
        RECT 28.085 200.025 28.870 200.195 ;
        RECT 29.145 199.745 29.355 200.275 ;
        RECT 29.620 199.960 29.950 200.485 ;
        RECT 30.460 200.400 30.860 200.485 ;
        RECT 31.525 200.985 31.795 201.375 ;
        RECT 31.985 201.155 32.200 202.295 ;
        RECT 32.370 201.155 32.705 202.125 ;
        RECT 32.875 201.990 33.125 202.295 ;
        RECT 35.880 202.275 45.540 202.445 ;
        RECT 32.875 201.650 34.030 201.990 ;
        RECT 32.875 201.155 33.125 201.650 ;
        RECT 36.055 201.605 36.225 202.105 ;
        RECT 36.395 201.775 36.725 202.275 ;
        RECT 36.055 201.435 36.720 201.605 ;
        RECT 31.525 200.655 32.320 200.985 ;
        RECT 30.120 199.745 30.290 200.355 ;
        RECT 30.460 199.965 30.790 200.400 ;
        RECT 31.525 200.275 31.725 200.655 ;
        RECT 32.490 200.545 32.705 201.155 ;
        RECT 35.970 200.615 36.320 201.265 ;
        RECT 30.960 199.745 31.130 200.260 ;
        RECT 31.465 200.005 31.725 200.275 ;
        RECT 31.950 199.745 32.280 200.485 ;
        RECT 32.450 199.925 32.705 200.545 ;
        RECT 32.875 200.330 33.125 200.565 ;
        RECT 36.490 200.445 36.720 201.435 ;
        RECT 32.875 200.020 34.030 200.330 ;
        RECT 36.055 200.275 36.720 200.445 ;
        RECT 32.875 199.745 33.125 200.020 ;
        RECT 36.055 199.985 36.225 200.275 ;
        RECT 11.140 199.575 20.800 199.745 ;
        RECT 23.560 199.575 33.220 199.745 ;
        RECT 36.395 199.725 36.725 200.105 ;
        RECT 36.895 199.985 37.080 202.105 ;
        RECT 37.320 201.815 37.585 202.275 ;
        RECT 37.755 201.680 38.005 202.105 ;
        RECT 38.215 201.830 39.320 202.000 ;
        RECT 37.700 201.550 38.005 201.680 ;
        RECT 37.250 200.355 37.530 201.305 ;
        RECT 37.700 200.445 37.870 201.550 ;
        RECT 38.040 200.765 38.280 201.360 ;
        RECT 38.450 201.295 38.980 201.660 ;
        RECT 38.450 200.595 38.620 201.295 ;
        RECT 39.150 201.215 39.320 201.830 ;
        RECT 39.490 201.475 39.660 202.275 ;
        RECT 39.830 201.775 40.080 202.105 ;
        RECT 40.305 201.805 41.190 201.975 ;
        RECT 39.150 201.125 39.660 201.215 ;
        RECT 37.700 200.315 37.925 200.445 ;
        RECT 38.095 200.375 38.620 200.595 ;
        RECT 38.790 200.955 39.660 201.125 ;
        RECT 37.335 199.725 37.585 200.185 ;
        RECT 37.755 200.175 37.925 200.315 ;
        RECT 38.790 200.175 38.960 200.955 ;
        RECT 39.490 200.885 39.660 200.955 ;
        RECT 39.170 200.705 39.370 200.735 ;
        RECT 39.830 200.705 40.000 201.775 ;
        RECT 40.170 200.885 40.360 201.605 ;
        RECT 39.170 200.405 40.000 200.705 ;
        RECT 40.530 200.675 40.850 201.635 ;
        RECT 37.755 200.005 38.090 200.175 ;
        RECT 38.285 200.005 38.960 200.175 ;
        RECT 39.280 199.725 39.650 200.225 ;
        RECT 39.830 200.175 40.000 200.405 ;
        RECT 40.385 200.345 40.850 200.675 ;
        RECT 41.020 200.965 41.190 201.805 ;
        RECT 41.370 201.775 41.685 202.275 ;
        RECT 41.920 201.545 42.260 202.105 ;
        RECT 41.360 201.170 42.260 201.545 ;
        RECT 42.430 201.265 42.600 202.275 ;
        RECT 42.070 200.965 42.260 201.170 ;
        RECT 42.770 201.215 43.100 202.060 ;
        RECT 43.270 201.360 43.445 202.275 ;
        RECT 43.785 201.355 44.115 202.085 ;
        RECT 42.770 201.135 43.180 201.215 ;
        RECT 42.945 201.085 43.180 201.135 ;
        RECT 41.020 200.635 41.900 200.965 ;
        RECT 42.070 200.635 42.820 200.965 ;
        RECT 41.020 200.175 41.190 200.635 ;
        RECT 42.070 200.465 42.270 200.635 ;
        RECT 42.990 200.505 43.180 201.085 ;
        RECT 42.935 200.465 43.180 200.505 ;
        RECT 39.830 200.005 40.235 200.175 ;
        RECT 40.405 200.005 41.190 200.175 ;
        RECT 41.465 199.725 41.675 200.255 ;
        RECT 41.940 199.940 42.270 200.465 ;
        RECT 42.780 200.380 43.180 200.465 ;
        RECT 43.845 200.965 44.115 201.355 ;
        RECT 44.305 201.135 44.520 202.275 ;
        RECT 44.690 201.135 45.025 202.105 ;
        RECT 45.195 202.010 45.445 202.275 ;
        RECT 45.195 201.570 46.690 202.010 ;
        RECT 45.195 201.135 45.445 201.570 ;
        RECT 133.285 201.325 133.455 203.230 ;
        RECT 134.515 203.060 134.775 203.230 ;
        RECT 135.025 203.110 135.325 203.570 ;
        RECT 136.005 203.390 136.175 205.205 ;
        RECT 133.730 202.890 134.775 203.060 ;
        RECT 134.995 202.910 135.325 203.110 ;
        RECT 135.505 203.020 136.175 203.390 ;
        RECT 133.730 201.955 133.900 202.890 ;
        RECT 134.070 202.360 134.435 202.720 ;
        RECT 134.605 202.700 134.775 202.890 ;
        RECT 134.605 202.530 135.725 202.700 ;
        RECT 134.070 202.190 135.355 202.360 ;
        RECT 134.370 201.780 134.965 202.020 ;
        RECT 135.135 201.835 135.355 202.190 ;
        RECT 135.555 202.025 135.725 202.530 ;
        RECT 133.625 201.610 134.180 201.745 ;
        RECT 135.555 201.665 135.725 201.830 ;
        RECT 135.285 201.610 135.725 201.665 ;
        RECT 133.625 201.495 135.725 201.610 ;
        RECT 134.050 201.440 135.415 201.495 ;
        RECT 136.005 201.325 136.175 203.020 ;
        RECT 43.845 200.635 44.640 200.965 ;
        RECT 42.440 199.725 42.610 200.335 ;
        RECT 42.780 199.945 43.110 200.380 ;
        RECT 43.845 200.255 44.045 200.635 ;
        RECT 44.810 200.525 45.025 201.135 ;
        RECT 133.285 201.060 133.915 201.325 ;
        RECT 43.280 199.725 43.450 200.240 ;
        RECT 43.785 199.985 44.045 200.255 ;
        RECT 44.270 199.725 44.600 200.465 ;
        RECT 44.770 199.905 45.025 200.525 ;
        RECT 45.195 200.380 45.445 200.545 ;
        RECT 133.285 200.465 133.455 201.060 ;
        RECT 134.425 200.990 135.375 201.270 ;
        RECT 135.545 201.075 136.175 201.325 ;
        RECT 133.625 200.635 135.745 200.820 ;
        RECT 136.005 200.465 136.175 201.075 ;
        RECT 45.195 200.010 46.100 200.380 ;
        RECT 133.285 200.135 133.955 200.465 ;
        RECT 134.125 200.230 135.455 200.460 ;
        RECT 45.195 199.725 45.445 200.010 ;
        RECT 35.880 199.555 45.540 199.725 ;
        RECT 133.285 199.535 133.455 200.135 ;
        RECT 134.125 199.965 134.295 200.230 ;
        RECT 133.625 199.795 134.295 199.965 ;
        RECT 134.465 199.710 135.115 200.060 ;
        RECT 135.285 199.965 135.455 200.230 ;
        RECT 135.625 200.135 136.175 200.465 ;
        RECT 135.285 199.795 135.745 199.965 ;
        RECT 133.285 199.245 134.620 199.535 ;
        RECT 133.285 199.075 133.455 199.245 ;
        RECT 133.285 198.825 134.595 199.075 ;
        RECT 133.285 198.150 133.455 198.825 ;
        RECT 134.810 198.660 134.990 199.710 ;
        RECT 136.005 199.535 136.175 200.135 ;
        RECT 135.280 199.245 136.175 199.535 ;
        RECT 136.005 199.075 136.175 199.245 ;
        RECT 135.185 198.825 136.175 199.075 ;
        RECT 134.740 198.655 134.990 198.660 ;
        RECT 133.625 198.440 135.825 198.655 ;
        RECT 133.625 198.320 134.595 198.440 ;
        RECT 135.205 198.400 135.825 198.440 ;
        RECT 133.285 197.935 134.595 198.150 ;
        RECT 133.285 197.075 133.455 197.935 ;
        RECT 134.765 197.745 135.095 198.270 ;
        RECT 136.005 198.230 136.175 198.825 ;
        RECT 135.265 197.900 136.175 198.230 ;
        RECT 133.645 197.675 135.095 197.745 ;
        RECT 133.645 197.475 135.745 197.675 ;
        RECT 133.645 197.415 134.375 197.475 ;
        RECT 135.475 197.415 135.745 197.475 ;
        RECT 136.005 197.080 136.175 197.900 ;
        RECT 133.285 196.900 134.370 197.075 ;
        RECT 135.490 196.910 136.175 197.080 ;
        RECT 96.530 196.550 96.880 196.570 ;
        RECT 96.530 196.545 97.090 196.550 ;
        RECT 96.530 196.375 108.070 196.545 ;
        RECT 96.530 196.370 97.090 196.375 ;
        RECT 96.530 195.600 96.880 196.370 ;
        RECT 97.310 195.185 97.480 196.375 ;
        RECT 97.650 195.820 97.950 196.205 ;
        RECT 98.120 195.995 98.450 196.375 ;
        RECT 99.000 195.945 99.340 196.375 ;
        RECT 97.650 195.275 98.040 195.820 ;
        RECT 99.510 195.775 99.735 196.205 ;
        RECT 100.015 195.995 100.360 196.375 ;
        RECT 100.540 195.825 100.710 196.115 ;
        RECT 100.880 195.915 101.130 196.375 ;
        RECT 98.235 195.605 99.735 195.775 ;
        RECT 96.420 193.870 96.940 194.610 ;
        RECT 97.310 193.870 97.480 194.670 ;
        RECT 97.650 194.565 97.820 195.275 ;
        RECT 98.235 195.065 98.405 195.605 ;
        RECT 99.080 195.535 99.735 195.605 ;
        RECT 99.910 195.655 100.710 195.825 ;
        RECT 101.300 195.865 102.170 196.205 ;
        RECT 97.990 194.735 98.405 195.065 ;
        RECT 97.650 194.050 98.030 194.565 ;
        RECT 96.420 193.825 97.480 193.870 ;
        RECT 98.200 193.825 98.370 194.565 ;
        RECT 98.575 194.005 98.910 195.435 ;
        RECT 99.080 194.625 99.250 195.535 ;
        RECT 99.910 195.065 100.080 195.655 ;
        RECT 101.300 195.485 101.470 195.865 ;
        RECT 102.405 195.745 102.575 196.205 ;
        RECT 102.745 195.915 103.115 196.375 ;
        RECT 103.410 195.775 103.580 196.115 ;
        RECT 103.750 195.945 104.080 196.375 ;
        RECT 104.315 195.775 104.485 196.115 ;
        RECT 100.250 195.315 101.470 195.485 ;
        RECT 101.640 195.405 102.100 195.695 ;
        RECT 102.405 195.575 102.965 195.745 ;
        RECT 103.410 195.605 104.485 195.775 ;
        RECT 104.655 195.875 105.335 196.205 ;
        RECT 105.550 195.875 105.800 196.205 ;
        RECT 105.970 195.915 106.220 196.375 ;
        RECT 106.420 196.190 106.680 196.375 ;
        RECT 102.795 195.435 102.965 195.575 ;
        RECT 101.640 195.395 102.605 195.405 ;
        RECT 101.300 195.225 101.470 195.315 ;
        RECT 101.930 195.235 102.605 195.395 ;
        RECT 99.420 195.035 100.080 195.065 ;
        RECT 99.420 194.815 100.255 195.035 ;
        RECT 99.910 194.735 100.255 194.815 ;
        RECT 99.080 194.455 99.735 194.625 ;
        RECT 99.080 193.825 99.315 194.285 ;
        RECT 99.485 194.085 99.735 194.455 ;
        RECT 100.085 194.205 100.255 194.735 ;
        RECT 100.425 194.775 100.965 195.145 ;
        RECT 101.300 195.055 101.705 195.225 ;
        RECT 100.425 194.375 100.665 194.775 ;
        RECT 101.145 194.605 101.365 194.885 ;
        RECT 100.835 194.435 101.365 194.605 ;
        RECT 100.835 194.205 101.005 194.435 ;
        RECT 101.535 194.275 101.705 195.055 ;
        RECT 101.875 194.445 102.225 195.065 ;
        RECT 102.395 194.445 102.605 195.235 ;
        RECT 102.795 195.265 104.295 195.435 ;
        RECT 102.795 194.575 102.965 195.265 ;
        RECT 104.655 195.095 104.825 195.875 ;
        RECT 105.630 195.745 105.800 195.875 ;
        RECT 103.135 194.925 104.825 195.095 ;
        RECT 104.995 195.315 105.460 195.705 ;
        RECT 105.630 195.575 106.025 195.745 ;
        RECT 103.135 194.745 103.305 194.925 ;
        RECT 100.085 194.035 101.005 194.205 ;
        RECT 101.175 193.825 101.365 194.265 ;
        RECT 101.535 193.995 102.485 194.275 ;
        RECT 102.795 194.185 103.055 194.575 ;
        RECT 103.475 194.505 104.265 194.755 ;
        RECT 102.705 194.015 103.055 194.185 ;
        RECT 103.265 193.825 103.595 194.285 ;
        RECT 104.470 194.215 104.640 194.925 ;
        RECT 104.995 194.725 105.165 195.315 ;
        RECT 104.810 194.505 105.165 194.725 ;
        RECT 105.335 194.505 105.685 195.125 ;
        RECT 105.855 194.215 106.025 195.575 ;
        RECT 106.390 195.405 106.715 196.190 ;
        RECT 106.195 194.355 106.655 195.405 ;
        RECT 104.470 194.045 105.325 194.215 ;
        RECT 105.530 194.045 106.025 194.215 ;
        RECT 106.195 193.825 106.525 194.185 ;
        RECT 106.885 194.085 107.055 196.205 ;
        RECT 107.225 195.875 107.555 196.375 ;
        RECT 133.285 196.230 133.455 196.900 ;
        RECT 134.515 196.740 135.350 196.810 ;
        RECT 134.515 196.730 135.785 196.740 ;
        RECT 133.670 196.620 135.785 196.730 ;
        RECT 133.670 196.575 134.645 196.620 ;
        RECT 133.670 196.400 134.595 196.575 ;
        RECT 135.225 196.565 135.785 196.620 ;
        RECT 107.725 195.705 107.980 196.205 ;
        RECT 107.230 195.535 107.980 195.705 ;
        RECT 133.285 196.060 134.465 196.230 ;
        RECT 107.230 194.545 107.460 195.535 ;
        RECT 107.630 195.350 107.980 195.365 ;
        RECT 107.630 194.750 110.570 195.350 ;
        RECT 133.285 195.315 133.455 196.060 ;
        RECT 134.765 195.900 135.095 196.450 ;
        RECT 135.265 196.410 135.785 196.565 ;
        RECT 136.005 196.240 136.175 196.910 ;
        RECT 135.395 196.070 136.175 196.240 ;
        RECT 134.765 195.890 135.790 195.900 ;
        RECT 133.625 195.700 135.790 195.890 ;
        RECT 133.625 195.550 134.560 195.700 ;
        RECT 135.265 195.570 135.790 195.700 ;
        RECT 133.285 195.000 133.955 195.315 ;
        RECT 107.630 194.715 107.980 194.750 ;
        RECT 107.230 194.375 107.980 194.545 ;
        RECT 107.225 193.825 107.555 194.205 ;
        RECT 107.725 194.085 107.980 194.375 ;
        RECT 96.420 193.655 108.070 193.825 ;
        RECT 96.420 193.640 97.330 193.655 ;
        RECT 133.285 193.290 133.455 195.000 ;
        RECT 134.185 194.990 134.560 195.550 ;
        RECT 134.765 194.820 135.095 195.530 ;
        RECT 136.005 195.305 136.175 196.070 ;
        RECT 135.475 195.095 136.175 195.305 ;
        RECT 133.755 194.650 135.725 194.820 ;
        RECT 133.755 193.935 133.925 194.650 ;
        RECT 134.095 194.160 135.385 194.480 ;
        RECT 135.055 194.015 135.385 194.160 ;
        RECT 135.555 194.035 135.725 194.650 ;
        RECT 134.125 193.800 134.845 193.990 ;
        RECT 133.625 193.630 133.955 193.710 ;
        RECT 135.555 193.630 135.725 193.865 ;
        RECT 133.625 193.460 135.725 193.630 ;
        RECT 133.285 193.120 134.255 193.290 ;
        RECT 134.515 193.120 134.845 193.290 ;
        RECT 98.070 192.195 98.830 192.220 ;
        RECT 98.070 192.025 101.530 192.195 ;
        RECT 98.070 192.000 98.830 192.025 ;
        RECT 98.070 191.550 98.440 192.000 ;
        RECT 99.055 191.355 99.335 192.025 ;
        RECT 98.855 190.730 99.170 191.155 ;
        RECT 99.505 191.135 99.805 191.685 ;
        RECT 100.015 191.305 100.345 192.025 ;
        RECT 100.535 191.305 100.985 191.855 ;
        RECT 99.505 190.965 100.445 191.135 ;
        RECT 98.855 190.715 99.320 190.730 ;
        RECT 100.275 190.715 100.445 190.965 ;
        RECT 98.855 190.465 99.545 190.715 ;
        RECT 99.775 190.465 100.105 190.715 ;
        RECT 100.275 190.385 100.565 190.715 ;
        RECT 100.735 190.670 100.985 191.305 ;
        RECT 101.155 190.885 101.445 192.025 ;
        RECT 103.390 192.005 105.690 192.175 ;
        RECT 103.520 190.865 103.785 192.005 ;
        RECT 103.955 191.035 104.285 191.835 ;
        RECT 104.455 191.205 104.625 192.005 ;
        RECT 104.795 191.055 105.125 191.835 ;
        RECT 105.295 191.545 105.505 192.005 ;
        RECT 133.285 191.215 133.455 193.120 ;
        RECT 134.515 192.950 134.775 193.120 ;
        RECT 135.025 193.000 135.325 193.460 ;
        RECT 136.005 193.280 136.175 195.095 ;
        RECT 133.730 192.780 134.775 192.950 ;
        RECT 134.995 192.800 135.325 193.000 ;
        RECT 135.505 192.910 136.175 193.280 ;
        RECT 133.730 191.845 133.900 192.780 ;
        RECT 134.070 192.250 134.435 192.610 ;
        RECT 134.605 192.590 134.775 192.780 ;
        RECT 134.605 192.420 135.725 192.590 ;
        RECT 134.070 192.080 135.355 192.250 ;
        RECT 134.370 191.670 134.965 191.910 ;
        RECT 135.135 191.725 135.355 192.080 ;
        RECT 135.555 191.915 135.725 192.420 ;
        RECT 133.625 191.500 134.180 191.635 ;
        RECT 135.555 191.555 135.725 191.720 ;
        RECT 135.285 191.500 135.725 191.555 ;
        RECT 133.625 191.385 135.725 191.500 ;
        RECT 134.050 191.330 135.415 191.385 ;
        RECT 136.005 191.215 136.175 192.910 ;
        RECT 104.795 191.035 105.560 191.055 ;
        RECT 103.955 190.865 105.560 191.035 ;
        RECT 103.495 190.670 105.125 190.695 ;
        RECT 100.735 190.450 105.125 190.670 ;
        RECT 98.240 189.480 98.780 190.300 ;
        RECT 100.275 190.295 100.445 190.385 ;
        RECT 99.055 190.105 100.445 190.295 ;
        RECT 99.055 189.745 99.385 190.105 ;
        RECT 100.735 189.935 100.985 190.450 ;
        RECT 103.495 190.445 105.125 190.450 ;
        RECT 105.295 190.275 105.560 190.865 ;
        RECT 98.240 189.475 98.980 189.480 ;
        RECT 100.015 189.475 100.265 189.935 ;
        RECT 100.435 189.645 100.985 189.935 ;
        RECT 101.155 189.475 101.445 190.275 ;
        RECT 103.955 190.095 105.560 190.275 ;
        RECT 133.285 190.950 133.915 191.215 ;
        RECT 133.285 190.355 133.455 190.950 ;
        RECT 134.425 190.880 135.375 191.160 ;
        RECT 135.545 190.965 136.175 191.215 ;
        RECT 133.625 190.525 135.745 190.710 ;
        RECT 136.005 190.355 136.175 190.965 ;
        RECT 98.240 189.305 101.530 189.475 ;
        RECT 103.520 189.455 103.785 189.915 ;
        RECT 103.955 189.625 104.285 190.095 ;
        RECT 104.455 189.455 104.625 189.915 ;
        RECT 104.795 189.625 105.125 190.095 ;
        RECT 133.285 190.025 133.955 190.355 ;
        RECT 134.125 190.120 135.455 190.350 ;
        RECT 105.295 189.455 105.545 189.920 ;
        RECT 133.285 189.510 133.455 190.025 ;
        RECT 134.125 189.855 134.295 190.120 ;
        RECT 133.625 189.685 134.295 189.855 ;
        RECT 134.465 189.600 135.115 189.950 ;
        RECT 135.285 189.855 135.455 190.120 ;
        RECT 135.625 190.025 136.175 190.355 ;
        RECT 135.285 189.685 135.745 189.855 ;
        RECT 136.005 189.650 136.175 190.025 ;
        RECT 98.240 189.300 98.980 189.305 ;
        RECT 103.390 189.285 105.690 189.455 ;
        RECT 134.580 188.230 135.080 189.600 ;
        RECT 136.005 189.510 136.200 189.650 ;
        RECT 136.010 189.340 136.200 189.510 ;
        RECT 135.390 188.820 136.200 189.340 ;
        RECT 96.270 187.795 96.990 187.820 ;
        RECT 96.270 187.625 107.950 187.795 ;
        RECT 96.270 187.590 96.990 187.625 ;
        RECT 96.290 186.710 96.700 187.590 ;
        RECT 97.190 186.435 97.360 187.625 ;
        RECT 97.530 187.070 97.830 187.455 ;
        RECT 98.000 187.245 98.330 187.625 ;
        RECT 98.880 187.195 99.220 187.625 ;
        RECT 97.530 186.525 97.920 187.070 ;
        RECT 99.390 187.025 99.615 187.455 ;
        RECT 99.895 187.245 100.240 187.625 ;
        RECT 100.420 187.075 100.590 187.365 ;
        RECT 100.760 187.165 101.010 187.625 ;
        RECT 98.115 186.855 99.615 187.025 ;
        RECT 96.330 185.090 96.730 185.790 ;
        RECT 97.190 185.090 97.360 185.920 ;
        RECT 97.530 185.815 97.700 186.525 ;
        RECT 98.115 186.315 98.285 186.855 ;
        RECT 98.960 186.785 99.615 186.855 ;
        RECT 99.790 186.905 100.590 187.075 ;
        RECT 101.180 187.115 102.050 187.455 ;
        RECT 97.870 185.985 98.285 186.315 ;
        RECT 97.530 185.300 97.910 185.815 ;
        RECT 96.310 185.075 97.360 185.090 ;
        RECT 98.080 185.075 98.250 185.815 ;
        RECT 98.455 185.255 98.790 186.685 ;
        RECT 98.960 185.875 99.130 186.785 ;
        RECT 99.790 186.315 99.960 186.905 ;
        RECT 101.180 186.735 101.350 187.115 ;
        RECT 102.285 186.995 102.455 187.455 ;
        RECT 102.625 187.165 102.995 187.625 ;
        RECT 103.290 187.025 103.460 187.365 ;
        RECT 103.630 187.195 103.960 187.625 ;
        RECT 104.195 187.025 104.365 187.365 ;
        RECT 100.130 186.565 101.350 186.735 ;
        RECT 101.520 186.655 101.980 186.945 ;
        RECT 102.285 186.825 102.845 186.995 ;
        RECT 103.290 186.855 104.365 187.025 ;
        RECT 104.535 187.125 105.215 187.455 ;
        RECT 105.430 187.125 105.680 187.455 ;
        RECT 105.850 187.165 106.100 187.625 ;
        RECT 106.310 187.440 106.570 187.625 ;
        RECT 102.675 186.685 102.845 186.825 ;
        RECT 101.520 186.645 102.485 186.655 ;
        RECT 101.180 186.475 101.350 186.565 ;
        RECT 101.810 186.485 102.485 186.645 ;
        RECT 99.300 186.285 99.960 186.315 ;
        RECT 99.300 186.065 100.135 186.285 ;
        RECT 99.790 185.985 100.135 186.065 ;
        RECT 98.960 185.705 99.615 185.875 ;
        RECT 98.960 185.075 99.195 185.535 ;
        RECT 99.365 185.335 99.615 185.705 ;
        RECT 99.965 185.455 100.135 185.985 ;
        RECT 100.305 186.025 100.845 186.395 ;
        RECT 101.180 186.305 101.585 186.475 ;
        RECT 100.305 185.625 100.545 186.025 ;
        RECT 101.025 185.855 101.245 186.135 ;
        RECT 100.715 185.685 101.245 185.855 ;
        RECT 100.715 185.455 100.885 185.685 ;
        RECT 101.415 185.525 101.585 186.305 ;
        RECT 101.755 185.695 102.105 186.315 ;
        RECT 102.275 185.695 102.485 186.485 ;
        RECT 102.675 186.515 104.175 186.685 ;
        RECT 102.675 185.825 102.845 186.515 ;
        RECT 104.535 186.345 104.705 187.125 ;
        RECT 105.510 186.995 105.680 187.125 ;
        RECT 103.015 186.175 104.705 186.345 ;
        RECT 104.875 186.565 105.340 186.955 ;
        RECT 105.510 186.825 105.905 186.995 ;
        RECT 103.015 185.995 103.185 186.175 ;
        RECT 99.965 185.285 100.885 185.455 ;
        RECT 101.055 185.075 101.245 185.515 ;
        RECT 101.415 185.245 102.365 185.525 ;
        RECT 102.675 185.435 102.935 185.825 ;
        RECT 103.355 185.755 104.145 186.005 ;
        RECT 102.585 185.265 102.935 185.435 ;
        RECT 103.145 185.075 103.475 185.535 ;
        RECT 104.350 185.465 104.520 186.175 ;
        RECT 104.875 185.975 105.045 186.565 ;
        RECT 104.690 185.755 105.045 185.975 ;
        RECT 105.215 185.755 105.565 186.375 ;
        RECT 105.735 185.465 105.905 186.825 ;
        RECT 106.270 186.655 106.595 187.440 ;
        RECT 106.075 185.605 106.535 186.655 ;
        RECT 104.350 185.295 105.205 185.465 ;
        RECT 105.410 185.295 105.905 185.465 ;
        RECT 106.075 185.075 106.405 185.435 ;
        RECT 106.765 185.335 106.935 187.455 ;
        RECT 107.105 187.125 107.435 187.625 ;
        RECT 107.605 186.955 107.860 187.455 ;
        RECT 107.110 186.785 107.860 186.955 ;
        RECT 107.110 185.795 107.340 186.785 ;
        RECT 107.510 186.610 107.860 186.615 ;
        RECT 107.510 185.980 110.450 186.610 ;
        RECT 107.510 185.970 109.740 185.980 ;
        RECT 107.510 185.965 107.860 185.970 ;
        RECT 107.110 185.625 107.860 185.795 ;
        RECT 107.105 185.075 107.435 185.455 ;
        RECT 107.605 185.335 107.860 185.625 ;
        RECT 96.310 184.905 107.950 185.075 ;
        RECT 96.310 184.900 97.280 184.905 ;
        RECT 87.440 150.400 97.940 150.450 ;
        RECT 87.390 150.280 97.940 150.400 ;
        RECT 87.390 150.120 97.980 150.280 ;
        RECT 98.450 150.200 104.570 150.440 ;
        RECT 78.580 150.000 85.070 150.010 ;
        RECT 78.580 149.980 86.110 150.000 ;
        RECT 68.990 149.975 69.560 149.980 ;
        RECT 58.090 149.810 69.560 149.975 ;
        RECT 58.090 149.805 69.130 149.810 ;
        RECT 53.690 148.780 55.780 149.320 ;
        RECT 58.180 149.135 58.435 149.635 ;
        RECT 58.605 149.305 58.935 149.805 ;
        RECT 58.180 148.965 58.930 149.135 ;
        RECT 58.180 148.780 58.530 148.795 ;
        RECT 53.690 148.170 58.530 148.780 ;
        RECT 53.690 147.220 55.780 148.170 ;
        RECT 58.180 148.145 58.530 148.170 ;
        RECT 58.700 147.975 58.930 148.965 ;
        RECT 58.180 147.805 58.930 147.975 ;
        RECT 58.180 147.515 58.435 147.805 ;
        RECT 58.605 147.255 58.935 147.635 ;
        RECT 59.105 147.515 59.275 149.635 ;
        RECT 59.450 149.620 59.770 149.805 ;
        RECT 59.445 148.835 59.770 149.620 ;
        RECT 59.940 149.345 60.190 149.805 ;
        RECT 60.360 149.305 60.610 149.635 ;
        RECT 60.825 149.305 61.505 149.635 ;
        RECT 60.360 149.175 60.530 149.305 ;
        RECT 60.135 149.005 60.530 149.175 ;
        RECT 59.505 147.785 59.965 148.835 ;
        RECT 60.135 147.645 60.305 149.005 ;
        RECT 60.700 148.745 61.165 149.135 ;
        RECT 60.475 147.935 60.825 148.555 ;
        RECT 60.995 148.155 61.165 148.745 ;
        RECT 61.335 148.525 61.505 149.305 ;
        RECT 61.675 149.205 61.845 149.545 ;
        RECT 62.080 149.375 62.410 149.805 ;
        RECT 62.580 149.205 62.750 149.545 ;
        RECT 63.045 149.345 63.415 149.805 ;
        RECT 61.675 149.035 62.750 149.205 ;
        RECT 63.585 149.175 63.755 149.635 ;
        RECT 63.990 149.295 64.860 149.635 ;
        RECT 65.030 149.345 65.280 149.805 ;
        RECT 63.195 149.005 63.755 149.175 ;
        RECT 63.195 148.865 63.365 149.005 ;
        RECT 61.865 148.695 63.365 148.865 ;
        RECT 64.060 148.835 64.520 149.125 ;
        RECT 61.335 148.355 63.025 148.525 ;
        RECT 60.995 147.935 61.350 148.155 ;
        RECT 61.520 147.645 61.690 148.355 ;
        RECT 61.895 147.935 62.685 148.185 ;
        RECT 62.855 148.175 63.025 148.355 ;
        RECT 63.195 148.005 63.365 148.695 ;
        RECT 59.635 147.255 59.965 147.615 ;
        RECT 60.135 147.475 60.630 147.645 ;
        RECT 60.835 147.475 61.690 147.645 ;
        RECT 62.565 147.255 62.895 147.715 ;
        RECT 63.105 147.615 63.365 148.005 ;
        RECT 63.555 148.825 64.520 148.835 ;
        RECT 64.690 148.915 64.860 149.295 ;
        RECT 65.450 149.255 65.620 149.545 ;
        RECT 65.800 149.425 66.145 149.805 ;
        RECT 65.450 149.085 66.250 149.255 ;
        RECT 63.555 148.665 64.230 148.825 ;
        RECT 64.690 148.745 65.910 148.915 ;
        RECT 63.555 147.875 63.765 148.665 ;
        RECT 64.690 148.655 64.860 148.745 ;
        RECT 63.935 147.875 64.285 148.495 ;
        RECT 64.455 148.485 64.860 148.655 ;
        RECT 64.455 147.705 64.625 148.485 ;
        RECT 64.795 148.035 65.015 148.315 ;
        RECT 65.195 148.205 65.735 148.575 ;
        RECT 66.080 148.495 66.250 149.085 ;
        RECT 66.425 149.205 66.650 149.635 ;
        RECT 66.820 149.375 67.160 149.805 ;
        RECT 67.710 149.425 68.040 149.805 ;
        RECT 68.210 149.250 68.510 149.635 ;
        RECT 66.425 149.035 67.925 149.205 ;
        RECT 66.425 148.965 67.080 149.035 ;
        RECT 66.080 148.465 66.740 148.495 ;
        RECT 64.795 147.865 65.325 148.035 ;
        RECT 63.105 147.445 63.455 147.615 ;
        RECT 63.675 147.425 64.625 147.705 ;
        RECT 64.795 147.255 64.985 147.695 ;
        RECT 65.155 147.635 65.325 147.865 ;
        RECT 65.495 147.805 65.735 148.205 ;
        RECT 65.905 148.245 66.740 148.465 ;
        RECT 65.905 148.165 66.250 148.245 ;
        RECT 65.905 147.635 66.075 148.165 ;
        RECT 66.910 148.055 67.080 148.965 ;
        RECT 65.155 147.465 66.075 147.635 ;
        RECT 66.425 147.885 67.080 148.055 ;
        RECT 66.425 147.515 66.675 147.885 ;
        RECT 66.845 147.255 67.080 147.715 ;
        RECT 67.250 147.435 67.585 148.865 ;
        RECT 67.755 148.495 67.925 149.035 ;
        RECT 68.120 148.705 68.510 149.250 ;
        RECT 67.755 148.165 68.170 148.495 ;
        RECT 68.340 147.995 68.510 148.705 ;
        RECT 68.680 148.615 68.850 149.805 ;
        RECT 69.385 149.230 69.555 149.810 ;
        RECT 72.760 149.805 75.520 149.975 ;
        RECT 78.580 149.840 86.120 149.980 ;
        RECT 87.390 149.860 88.360 150.120 ;
        RECT 70.990 148.500 71.940 148.800 ;
        RECT 72.890 148.665 73.155 149.805 ;
        RECT 73.325 148.835 73.655 149.635 ;
        RECT 73.825 149.005 73.995 149.805 ;
        RECT 74.165 148.855 74.495 149.635 ;
        RECT 74.665 149.345 74.875 149.805 ;
        RECT 74.165 148.835 74.930 148.855 ;
        RECT 73.325 148.665 74.930 148.835 ;
        RECT 70.970 148.490 71.940 148.500 ;
        RECT 72.865 148.490 74.495 148.495 ;
        RECT 70.970 148.245 74.495 148.490 ;
        RECT 74.665 148.455 74.930 148.665 ;
        RECT 75.145 148.640 75.435 149.805 ;
        RECT 75.710 148.455 76.330 148.550 ;
        RECT 70.970 148.240 73.180 148.245 ;
        RECT 70.990 148.230 73.180 148.240 ;
        RECT 67.790 147.255 67.960 147.995 ;
        RECT 68.130 147.480 68.510 147.995 ;
        RECT 68.680 147.255 68.850 148.100 ;
        RECT 69.210 148.010 70.130 148.160 ;
        RECT 70.990 148.120 71.940 148.230 ;
        RECT 74.665 148.155 76.330 148.455 ;
        RECT 74.665 148.075 74.930 148.155 ;
        RECT 69.190 147.520 70.130 148.010 ;
        RECT 73.325 147.895 74.930 148.075 ;
        RECT 69.210 147.510 70.130 147.520 ;
        RECT 72.890 147.255 73.155 147.715 ;
        RECT 73.325 147.425 73.655 147.895 ;
        RECT 73.825 147.255 73.995 147.715 ;
        RECT 74.165 147.425 74.495 147.895 ;
        RECT 74.665 147.255 74.915 147.720 ;
        RECT 75.145 147.255 75.435 147.980 ;
        RECT 75.710 147.930 76.330 148.155 ;
        RECT 58.090 147.085 69.130 147.255 ;
        RECT 72.760 147.085 75.520 147.255 ;
        RECT 78.580 146.350 78.750 149.840 ;
        RECT 79.290 149.330 79.620 149.500 ;
        RECT 79.150 147.075 79.320 149.115 ;
        RECT 79.590 148.210 79.760 149.115 ;
        RECT 80.160 148.210 80.330 149.840 ;
        RECT 80.870 149.330 81.200 149.500 ;
        RECT 80.730 148.210 80.900 149.115 ;
        RECT 79.590 147.970 80.900 148.210 ;
        RECT 79.590 147.075 79.760 147.970 ;
        RECT 79.290 146.690 79.620 146.860 ;
        RECT 80.160 146.350 80.330 147.970 ;
        RECT 80.730 147.075 80.900 147.970 ;
        RECT 81.170 147.075 81.340 149.115 ;
        RECT 81.740 148.190 81.910 149.840 ;
        RECT 82.450 149.330 82.780 149.500 ;
        RECT 82.310 148.190 82.480 149.115 ;
        RECT 81.730 147.960 82.480 148.190 ;
        RECT 80.870 146.690 81.200 146.860 ;
        RECT 81.740 146.350 81.910 147.960 ;
        RECT 82.310 147.075 82.480 147.960 ;
        RECT 82.750 147.075 82.920 149.115 ;
        RECT 82.450 146.690 82.780 146.860 ;
        RECT 83.320 146.350 83.490 149.840 ;
        RECT 84.900 149.670 86.120 149.840 ;
        RECT 84.900 149.650 86.110 149.670 ;
        RECT 84.030 149.330 84.360 149.500 ;
        RECT 83.890 147.075 84.060 149.115 ;
        RECT 84.330 147.075 84.500 149.115 ;
        RECT 84.030 146.690 84.360 146.860 ;
        RECT 84.900 146.350 85.070 149.650 ;
        RECT 87.380 149.610 88.360 149.860 ;
        RECT 88.580 150.110 90.330 150.120 ;
        RECT 88.580 149.610 88.750 150.110 ;
        RECT 87.380 149.300 88.750 149.610 ;
        RECT 89.290 149.600 89.620 149.770 ;
        RECT 87.380 148.980 88.760 149.300 ;
        RECT 87.380 148.970 88.340 148.980 ;
        RECT 67.170 146.275 68.490 146.310 ;
        RECT 60.260 146.055 62.560 146.225 ;
        RECT 64.970 146.105 68.490 146.275 ;
        RECT 78.580 146.180 85.070 146.350 ;
        RECT 87.400 147.290 88.130 148.970 ;
        RECT 88.580 147.820 88.750 148.980 ;
        RECT 89.150 148.545 89.320 149.385 ;
        RECT 89.590 149.070 89.760 149.385 ;
        RECT 90.160 149.070 90.330 150.110 ;
        RECT 89.590 148.830 90.330 149.070 ;
        RECT 89.590 148.545 89.760 148.830 ;
        RECT 89.290 148.160 89.620 148.330 ;
        RECT 90.160 147.820 90.330 148.830 ;
        RECT 88.580 147.650 90.330 147.820 ;
        RECT 90.690 150.100 92.440 150.120 ;
        RECT 90.690 147.810 90.860 150.100 ;
        RECT 91.400 149.590 91.730 149.760 ;
        RECT 91.260 148.535 91.430 149.375 ;
        RECT 91.700 149.040 91.870 149.375 ;
        RECT 92.270 149.040 92.440 150.100 ;
        RECT 91.700 148.800 92.440 149.040 ;
        RECT 91.700 148.535 91.870 148.800 ;
        RECT 91.400 148.150 91.730 148.320 ;
        RECT 92.270 147.810 92.440 148.800 ;
        RECT 90.690 147.640 92.440 147.810 ;
        RECT 92.800 150.110 94.550 150.120 ;
        RECT 92.800 147.820 92.970 150.110 ;
        RECT 93.510 149.600 93.840 149.770 ;
        RECT 93.370 148.545 93.540 149.385 ;
        RECT 93.810 149.030 93.980 149.385 ;
        RECT 94.380 149.030 94.550 150.110 ;
        RECT 93.800 148.790 94.550 149.030 ;
        RECT 93.810 148.545 93.980 148.790 ;
        RECT 93.510 148.160 93.840 148.330 ;
        RECT 94.380 147.820 94.550 148.790 ;
        RECT 92.800 147.650 94.550 147.820 ;
        RECT 96.230 150.110 97.980 150.120 ;
        RECT 96.230 149.090 96.400 150.110 ;
        RECT 96.940 149.600 97.270 149.770 ;
        RECT 96.800 149.090 96.970 149.385 ;
        RECT 96.230 148.850 96.970 149.090 ;
        RECT 96.230 147.820 96.400 148.850 ;
        RECT 96.800 148.545 96.970 148.850 ;
        RECT 97.240 148.545 97.410 149.385 ;
        RECT 96.940 148.160 97.270 148.330 ;
        RECT 97.810 147.820 97.980 150.110 ;
        RECT 96.230 147.650 97.980 147.820 ;
        RECT 98.370 149.980 104.570 150.200 ;
        RECT 98.370 147.830 98.540 149.980 ;
        RECT 99.170 149.520 101.170 149.690 ;
        RECT 98.940 148.510 99.110 149.350 ;
        RECT 101.230 149.040 101.400 149.350 ;
        RECT 101.800 149.040 101.970 149.980 ;
        RECT 101.230 148.800 101.970 149.040 ;
        RECT 103.610 148.960 104.570 149.980 ;
        RECT 101.230 148.510 101.400 148.800 ;
        RECT 99.170 148.170 101.170 148.340 ;
        RECT 101.800 147.830 101.970 148.800 ;
        RECT 98.370 147.660 101.970 147.830 ;
        RECT 87.400 147.120 99.780 147.290 ;
        RECT 60.445 145.595 60.655 146.055 ;
        RECT 60.825 145.105 61.155 145.885 ;
        RECT 61.325 145.255 61.495 146.055 ;
        RECT 60.390 145.085 61.155 145.105 ;
        RECT 61.665 145.085 61.995 145.885 ;
        RECT 59.230 144.940 59.960 144.970 ;
        RECT 60.390 144.940 61.995 145.085 ;
        RECT 59.230 144.915 61.995 144.940 ;
        RECT 62.165 144.915 62.430 146.055 ;
        RECT 65.055 144.965 65.345 146.105 ;
        RECT 65.515 145.385 65.965 145.935 ;
        RECT 66.155 145.385 66.485 146.105 ;
        RECT 67.165 146.100 68.490 146.105 ;
        RECT 59.230 144.350 60.655 144.915 ;
        RECT 63.940 144.790 64.780 144.800 ;
        RECT 65.515 144.790 65.765 145.385 ;
        RECT 66.695 145.215 66.995 145.765 ;
        RECT 67.165 145.435 67.445 146.100 ;
        RECT 68.120 146.070 68.490 146.100 ;
        RECT 68.120 145.900 68.510 146.070 ;
        RECT 68.335 145.320 68.505 145.900 ;
        RECT 87.400 145.720 88.130 147.120 ;
        RECT 88.460 146.250 88.630 146.580 ;
        RECT 88.845 146.550 98.885 146.720 ;
        RECT 88.845 146.110 98.885 146.280 ;
        RECT 99.100 146.250 99.270 146.580 ;
        RECT 87.400 145.710 88.180 145.720 ;
        RECT 99.610 145.710 99.780 147.120 ;
        RECT 103.630 145.960 104.510 146.070 ;
        RECT 78.580 145.520 85.670 145.690 ;
        RECT 66.055 145.045 66.995 145.215 ;
        RECT 67.330 145.120 67.645 145.235 ;
        RECT 71.090 145.120 72.140 145.390 ;
        RECT 66.055 144.795 66.225 145.045 ;
        RECT 66.410 144.795 66.750 144.860 ;
        RECT 67.330 144.795 72.140 145.120 ;
        RECT 60.825 144.740 62.455 144.745 ;
        RECT 63.940 144.740 65.765 144.790 ;
        RECT 60.825 144.530 65.765 144.740 ;
        RECT 60.825 144.520 64.880 144.530 ;
        RECT 60.825 144.495 64.780 144.520 ;
        RECT 62.110 144.490 64.780 144.495 ;
        RECT 63.940 144.480 64.780 144.490 ;
        RECT 59.230 144.300 59.960 144.350 ;
        RECT 60.390 144.325 60.655 144.350 ;
        RECT 60.390 144.145 61.995 144.325 ;
        RECT 60.405 143.505 60.655 143.970 ;
        RECT 60.825 143.675 61.155 144.145 ;
        RECT 61.325 143.505 61.495 143.965 ;
        RECT 61.665 143.675 61.995 144.145 ;
        RECT 62.165 143.505 62.430 143.965 ;
        RECT 65.055 143.555 65.345 144.355 ;
        RECT 65.515 144.015 65.765 144.530 ;
        RECT 65.935 144.465 66.225 144.795 ;
        RECT 66.395 144.550 66.750 144.795 ;
        RECT 66.955 144.560 72.140 144.795 ;
        RECT 66.395 144.545 66.725 144.550 ;
        RECT 66.955 144.545 67.645 144.560 ;
        RECT 71.090 144.500 72.140 144.560 ;
        RECT 66.055 144.375 66.225 144.465 ;
        RECT 66.055 144.185 67.445 144.375 ;
        RECT 65.515 143.725 66.065 144.015 ;
        RECT 66.235 143.555 66.485 144.015 ;
        RECT 67.115 143.825 67.445 144.185 ;
        RECT 67.890 143.820 68.730 144.370 ;
        RECT 78.580 144.320 78.750 145.520 ;
        RECT 79.365 145.010 79.695 145.180 ;
        RECT 79.150 144.320 79.320 144.840 ;
        RECT 78.580 144.110 79.320 144.320 ;
        RECT 60.260 143.335 62.560 143.505 ;
        RECT 64.970 143.385 67.730 143.555 ;
        RECT 78.580 143.120 78.750 144.110 ;
        RECT 79.150 143.800 79.320 144.110 ;
        RECT 79.740 143.800 79.910 144.840 ;
        RECT 80.310 144.320 80.480 145.520 ;
        RECT 81.095 145.010 81.425 145.180 ;
        RECT 80.880 144.320 81.050 144.840 ;
        RECT 80.310 144.110 81.050 144.320 ;
        RECT 79.365 143.460 79.695 143.630 ;
        RECT 80.310 143.120 80.480 144.110 ;
        RECT 80.880 143.800 81.050 144.110 ;
        RECT 81.470 143.800 81.640 144.840 ;
        RECT 82.040 144.310 82.210 145.520 ;
        RECT 82.825 145.010 83.155 145.180 ;
        RECT 82.610 144.310 82.780 144.840 ;
        RECT 82.040 144.100 82.780 144.310 ;
        RECT 81.095 143.460 81.425 143.630 ;
        RECT 82.040 143.120 82.210 144.100 ;
        RECT 82.610 143.800 82.780 144.100 ;
        RECT 83.200 143.800 83.370 144.840 ;
        RECT 82.825 143.460 83.155 143.630 ;
        RECT 83.770 143.120 83.940 145.520 ;
        RECT 84.555 145.010 84.885 145.180 ;
        RECT 84.340 143.800 84.510 144.840 ;
        RECT 84.930 143.800 85.100 144.840 ;
        RECT 84.555 143.460 84.885 143.630 ;
        RECT 85.500 143.270 85.670 145.520 ;
        RECT 87.400 145.540 99.780 145.710 ;
        RECT 100.150 145.790 104.510 145.960 ;
        RECT 85.500 143.120 86.470 143.270 ;
        RECT 78.580 142.950 86.470 143.120 ;
        RECT 87.400 143.050 88.180 145.540 ;
        RECT 93.050 145.010 99.790 145.180 ;
        RECT 93.050 143.600 93.220 145.010 ;
        RECT 93.560 144.140 93.730 144.470 ;
        RECT 93.900 144.440 98.940 144.610 ;
        RECT 93.900 144.000 98.940 144.170 ;
        RECT 99.110 144.140 99.280 144.470 ;
        RECT 99.620 143.600 99.790 145.010 ;
        RECT 93.050 143.430 99.790 143.600 ;
        RECT 100.150 143.590 100.320 145.790 ;
        RECT 100.950 145.280 102.950 145.450 ;
        RECT 100.720 144.270 100.890 145.110 ;
        RECT 103.010 145.070 103.180 145.110 ;
        RECT 103.580 145.070 104.510 145.790 ;
        RECT 103.010 144.280 104.510 145.070 ;
        RECT 103.010 144.270 103.180 144.280 ;
        RECT 100.950 143.930 102.950 144.100 ;
        RECT 103.580 143.770 104.510 144.280 ;
        RECT 103.580 143.590 103.750 143.770 ;
        RECT 100.150 143.420 103.750 143.590 ;
        RECT 87.400 142.920 99.770 143.050 ;
        RECT 87.420 142.880 99.770 142.920 ;
        RECT 87.420 142.870 88.180 142.880 ;
        RECT 68.440 142.565 69.480 142.580 ;
        RECT 57.860 142.395 69.480 142.565 ;
        RECT 57.950 141.725 58.205 142.225 ;
        RECT 58.375 141.895 58.705 142.395 ;
        RECT 57.950 141.555 58.700 141.725 ;
        RECT 54.260 141.380 55.090 141.390 ;
        RECT 57.950 141.380 58.300 141.385 ;
        RECT 54.260 141.370 58.300 141.380 ;
        RECT 53.880 140.740 58.300 141.370 ;
        RECT 53.880 138.310 55.640 140.740 ;
        RECT 57.950 140.735 58.300 140.740 ;
        RECT 58.470 140.565 58.700 141.555 ;
        RECT 57.950 140.395 58.700 140.565 ;
        RECT 57.950 140.105 58.205 140.395 ;
        RECT 58.375 139.845 58.705 140.225 ;
        RECT 58.875 140.105 59.045 142.225 ;
        RECT 59.220 142.210 59.530 142.395 ;
        RECT 59.215 141.425 59.540 142.210 ;
        RECT 59.710 141.935 59.960 142.395 ;
        RECT 60.130 141.895 60.380 142.225 ;
        RECT 60.595 141.895 61.275 142.225 ;
        RECT 60.130 141.765 60.300 141.895 ;
        RECT 59.905 141.595 60.300 141.765 ;
        RECT 59.275 140.375 59.735 141.425 ;
        RECT 59.905 140.235 60.075 141.595 ;
        RECT 60.470 141.335 60.935 141.725 ;
        RECT 60.245 140.525 60.595 141.145 ;
        RECT 60.765 140.745 60.935 141.335 ;
        RECT 61.105 141.115 61.275 141.895 ;
        RECT 61.445 141.795 61.615 142.135 ;
        RECT 61.850 141.965 62.180 142.395 ;
        RECT 62.350 141.795 62.520 142.135 ;
        RECT 62.815 141.935 63.185 142.395 ;
        RECT 61.445 141.625 62.520 141.795 ;
        RECT 63.355 141.765 63.525 142.225 ;
        RECT 63.760 141.885 64.630 142.225 ;
        RECT 64.800 141.935 65.050 142.395 ;
        RECT 62.965 141.595 63.525 141.765 ;
        RECT 62.965 141.455 63.135 141.595 ;
        RECT 61.635 141.285 63.135 141.455 ;
        RECT 63.830 141.425 64.290 141.715 ;
        RECT 61.105 140.945 62.795 141.115 ;
        RECT 60.765 140.525 61.120 140.745 ;
        RECT 61.290 140.235 61.460 140.945 ;
        RECT 61.665 140.525 62.455 140.775 ;
        RECT 62.625 140.765 62.795 140.945 ;
        RECT 62.965 140.595 63.135 141.285 ;
        RECT 59.405 139.845 59.735 140.205 ;
        RECT 59.905 140.065 60.400 140.235 ;
        RECT 60.605 140.065 61.460 140.235 ;
        RECT 62.335 139.845 62.665 140.305 ;
        RECT 62.875 140.205 63.135 140.595 ;
        RECT 63.325 141.415 64.290 141.425 ;
        RECT 64.460 141.505 64.630 141.885 ;
        RECT 65.220 141.845 65.390 142.135 ;
        RECT 65.570 142.015 65.915 142.395 ;
        RECT 65.220 141.675 66.020 141.845 ;
        RECT 63.325 141.255 64.000 141.415 ;
        RECT 64.460 141.335 65.680 141.505 ;
        RECT 63.325 140.465 63.535 141.255 ;
        RECT 64.460 141.245 64.630 141.335 ;
        RECT 63.705 140.465 64.055 141.085 ;
        RECT 64.225 141.075 64.630 141.245 ;
        RECT 64.225 140.295 64.395 141.075 ;
        RECT 64.565 140.625 64.785 140.905 ;
        RECT 64.965 140.795 65.505 141.165 ;
        RECT 65.850 141.085 66.020 141.675 ;
        RECT 66.195 141.795 66.420 142.225 ;
        RECT 66.590 141.965 66.930 142.395 ;
        RECT 67.480 142.015 67.810 142.395 ;
        RECT 68.440 142.390 69.480 142.395 ;
        RECT 67.980 141.840 68.280 142.225 ;
        RECT 66.195 141.625 67.695 141.795 ;
        RECT 66.195 141.555 66.850 141.625 ;
        RECT 65.850 141.055 66.510 141.085 ;
        RECT 64.565 140.455 65.095 140.625 ;
        RECT 62.875 140.035 63.225 140.205 ;
        RECT 63.445 140.015 64.395 140.295 ;
        RECT 64.565 139.845 64.755 140.285 ;
        RECT 64.925 140.225 65.095 140.455 ;
        RECT 65.265 140.395 65.505 140.795 ;
        RECT 65.675 140.835 66.510 141.055 ;
        RECT 65.675 140.755 66.020 140.835 ;
        RECT 65.675 140.225 65.845 140.755 ;
        RECT 66.680 140.645 66.850 141.555 ;
        RECT 64.925 140.055 65.845 140.225 ;
        RECT 66.195 140.475 66.850 140.645 ;
        RECT 66.195 140.105 66.445 140.475 ;
        RECT 66.615 139.845 66.850 140.305 ;
        RECT 67.020 140.025 67.355 141.455 ;
        RECT 67.525 141.085 67.695 141.625 ;
        RECT 67.890 141.295 68.280 141.840 ;
        RECT 67.525 140.755 67.940 141.085 ;
        RECT 68.110 140.585 68.280 141.295 ;
        RECT 68.450 141.205 68.620 142.390 ;
        RECT 69.070 142.360 69.470 142.390 ;
        RECT 69.295 141.780 69.465 142.360 ;
        RECT 87.420 141.490 88.130 142.870 ;
        RECT 88.450 142.010 88.620 142.340 ;
        RECT 88.835 142.310 98.875 142.480 ;
        RECT 88.835 141.870 98.875 142.040 ;
        RECT 99.090 142.010 99.260 142.340 ;
        RECT 87.420 141.470 88.180 141.490 ;
        RECT 99.600 141.470 99.770 142.880 ;
        RECT 87.420 141.300 99.770 141.470 ;
        RECT 100.130 141.640 103.730 141.720 ;
        RECT 100.130 141.550 104.530 141.640 ;
        RECT 67.560 139.845 67.730 140.585 ;
        RECT 67.900 140.070 68.280 140.585 ;
        RECT 68.450 139.845 68.620 140.690 ;
        RECT 69.220 140.640 69.870 140.820 ;
        RECT 57.860 139.675 68.900 139.845 ;
        RECT 69.200 139.730 69.880 140.640 ;
        RECT 87.420 138.820 88.180 141.300 ;
        RECT 93.030 140.900 99.770 140.930 ;
        RECT 100.130 140.900 100.300 141.550 ;
        RECT 100.930 141.040 102.930 141.210 ;
        RECT 93.030 140.760 100.300 140.900 ;
        RECT 93.030 139.350 93.200 140.760 ;
        RECT 93.540 139.890 93.710 140.220 ;
        RECT 93.880 140.190 98.920 140.360 ;
        RECT 93.880 139.750 98.920 139.920 ;
        RECT 99.090 139.890 99.260 140.220 ;
        RECT 99.600 139.350 100.300 140.760 ;
        RECT 100.700 140.030 100.870 140.870 ;
        RECT 102.990 140.830 103.160 140.870 ;
        RECT 103.560 140.830 104.530 141.550 ;
        RECT 102.990 140.040 104.530 140.830 ;
        RECT 102.990 140.030 103.160 140.040 ;
        RECT 100.930 139.690 102.930 139.860 ;
        RECT 103.560 139.350 104.530 140.040 ;
        RECT 93.030 139.340 104.530 139.350 ;
        RECT 93.030 139.200 103.730 139.340 ;
        RECT 93.030 139.180 99.770 139.200 ;
        RECT 100.130 139.180 103.730 139.200 ;
        RECT 87.420 138.650 99.770 138.820 ;
        RECT 87.420 138.640 88.180 138.650 ;
        RECT 87.420 138.630 88.160 138.640 ;
        RECT 71.120 138.605 71.530 138.610 ;
        RECT 71.120 138.525 81.090 138.605 ;
        RECT 70.400 138.435 81.090 138.525 ;
        RECT 70.400 138.355 71.775 138.435 ;
        RECT 53.900 138.300 55.630 138.310 ;
        RECT 70.400 137.565 70.570 138.355 ;
        RECT 71.120 138.340 71.775 138.355 ;
        RECT 70.400 137.395 71.245 137.565 ;
        RECT 71.525 137.295 71.775 138.340 ;
        RECT 71.945 137.295 72.280 138.265 ;
        RECT 72.450 137.295 72.665 138.435 ;
        RECT 72.855 137.515 73.185 138.245 ;
        RECT 73.525 137.520 73.700 138.435 ;
        RECT 70.920 135.890 71.290 136.730 ;
        RECT 71.525 135.890 71.775 136.705 ;
        RECT 71.945 136.685 72.160 137.295 ;
        RECT 72.855 137.125 73.125 137.515 ;
        RECT 73.870 137.375 74.200 138.220 ;
        RECT 74.370 137.425 74.540 138.435 ;
        RECT 74.710 137.705 75.050 138.265 ;
        RECT 75.285 137.935 75.600 138.435 ;
        RECT 75.780 137.965 76.665 138.135 ;
        RECT 72.330 136.795 73.125 137.125 ;
        RECT 71.945 136.065 72.200 136.685 ;
        RECT 70.920 135.885 71.775 135.890 ;
        RECT 72.370 135.885 72.700 136.625 ;
        RECT 72.925 136.415 73.125 136.795 ;
        RECT 73.790 137.295 74.200 137.375 ;
        RECT 74.710 137.330 75.610 137.705 ;
        RECT 73.790 137.245 74.025 137.295 ;
        RECT 73.790 136.665 73.980 137.245 ;
        RECT 74.710 137.125 74.900 137.330 ;
        RECT 75.780 137.125 75.950 137.965 ;
        RECT 76.890 137.935 77.140 138.265 ;
        RECT 74.150 136.795 74.900 137.125 ;
        RECT 75.070 136.795 75.950 137.125 ;
        RECT 73.790 136.625 74.035 136.665 ;
        RECT 74.700 136.625 74.900 136.795 ;
        RECT 73.790 136.540 74.190 136.625 ;
        RECT 72.925 136.145 73.185 136.415 ;
        RECT 73.520 135.885 73.690 136.400 ;
        RECT 73.860 136.105 74.190 136.540 ;
        RECT 74.360 135.885 74.530 136.495 ;
        RECT 74.700 136.100 75.030 136.625 ;
        RECT 75.295 135.885 75.505 136.415 ;
        RECT 75.780 136.335 75.950 136.795 ;
        RECT 76.120 136.835 76.440 137.795 ;
        RECT 76.610 137.045 76.800 137.765 ;
        RECT 76.970 136.865 77.140 137.935 ;
        RECT 77.310 137.635 77.480 138.435 ;
        RECT 77.650 137.990 78.755 138.160 ;
        RECT 77.650 137.375 77.820 137.990 ;
        RECT 78.965 137.840 79.215 138.265 ;
        RECT 79.385 137.975 79.650 138.435 ;
        RECT 77.990 137.455 78.520 137.820 ;
        RECT 78.965 137.710 79.270 137.840 ;
        RECT 77.310 137.285 77.820 137.375 ;
        RECT 77.310 137.115 78.180 137.285 ;
        RECT 77.310 137.045 77.480 137.115 ;
        RECT 77.600 136.865 77.800 136.895 ;
        RECT 76.120 136.505 76.585 136.835 ;
        RECT 76.970 136.565 77.800 136.865 ;
        RECT 76.970 136.335 77.140 136.565 ;
        RECT 75.780 136.165 76.565 136.335 ;
        RECT 76.735 136.165 77.140 136.335 ;
        RECT 77.320 135.885 77.690 136.385 ;
        RECT 78.010 136.335 78.180 137.115 ;
        RECT 78.350 136.755 78.520 137.455 ;
        RECT 78.690 136.925 78.930 137.520 ;
        RECT 78.350 136.535 78.875 136.755 ;
        RECT 79.100 136.605 79.270 137.710 ;
        RECT 79.045 136.475 79.270 136.605 ;
        RECT 79.440 136.515 79.720 137.465 ;
        RECT 79.045 136.335 79.215 136.475 ;
        RECT 78.010 136.165 78.685 136.335 ;
        RECT 78.880 136.165 79.215 136.335 ;
        RECT 79.385 135.885 79.635 136.345 ;
        RECT 79.890 136.145 80.075 138.265 ;
        RECT 80.245 137.935 80.575 138.435 ;
        RECT 80.745 137.765 80.915 138.265 ;
        RECT 80.250 137.595 80.915 137.765 ;
        RECT 80.250 136.605 80.480 137.595 ;
        RECT 80.650 137.070 81.000 137.425 ;
        RECT 87.430 137.280 88.160 138.630 ;
        RECT 88.450 137.780 88.620 138.110 ;
        RECT 88.835 138.080 98.875 138.250 ;
        RECT 88.835 137.640 98.875 137.810 ;
        RECT 99.090 137.780 99.260 138.110 ;
        RECT 87.430 137.240 90.050 137.280 ;
        RECT 99.600 137.240 99.770 138.650 ;
        RECT 87.430 137.070 99.770 137.240 ;
        RECT 100.140 137.310 104.490 137.480 ;
        RECT 80.650 136.890 82.690 137.070 ;
        RECT 80.650 136.775 81.000 136.890 ;
        RECT 87.430 136.790 90.050 137.070 ;
        RECT 80.250 136.435 80.915 136.605 ;
        RECT 80.245 135.890 80.575 136.265 ;
        RECT 80.745 136.145 80.915 136.435 ;
        RECT 89.870 136.565 90.050 136.790 ;
        RECT 89.870 136.370 91.185 136.565 ;
        RECT 89.875 136.335 91.185 136.370 ;
        RECT 80.245 135.885 81.550 135.890 ;
        RECT 70.920 135.720 81.550 135.885 ;
        RECT 71.430 135.715 81.090 135.720 ;
        RECT 71.050 135.085 71.510 135.090 ;
        RECT 71.050 134.990 81.070 135.085 ;
        RECT 69.865 134.920 81.070 134.990 ;
        RECT 69.865 134.820 71.220 134.920 ;
        RECT 71.410 134.915 81.070 134.920 ;
        RECT 69.865 134.030 70.035 134.820 ;
        RECT 69.865 133.860 70.710 134.030 ;
        RECT 71.505 133.775 71.755 134.915 ;
        RECT 71.925 133.775 72.260 134.745 ;
        RECT 72.430 133.775 72.645 134.915 ;
        RECT 72.835 133.995 73.165 134.725 ;
        RECT 73.505 134.000 73.680 134.915 ;
        RECT 70.920 132.480 71.270 133.250 ;
        RECT 71.505 132.480 71.755 133.185 ;
        RECT 71.925 133.165 72.140 133.775 ;
        RECT 72.835 133.605 73.105 133.995 ;
        RECT 73.850 133.855 74.180 134.700 ;
        RECT 74.350 133.905 74.520 134.915 ;
        RECT 74.690 134.185 75.030 134.745 ;
        RECT 75.265 134.415 75.580 134.915 ;
        RECT 75.760 134.445 76.645 134.615 ;
        RECT 72.310 133.275 73.105 133.605 ;
        RECT 71.925 132.545 72.180 133.165 ;
        RECT 70.930 132.365 71.755 132.480 ;
        RECT 72.350 132.365 72.680 133.105 ;
        RECT 72.905 132.895 73.105 133.275 ;
        RECT 73.770 133.775 74.180 133.855 ;
        RECT 74.690 133.810 75.590 134.185 ;
        RECT 73.770 133.725 74.005 133.775 ;
        RECT 73.770 133.145 73.960 133.725 ;
        RECT 74.690 133.605 74.880 133.810 ;
        RECT 75.760 133.605 75.930 134.445 ;
        RECT 76.870 134.415 77.120 134.745 ;
        RECT 74.130 133.275 74.880 133.605 ;
        RECT 75.050 133.275 75.930 133.605 ;
        RECT 73.770 133.105 74.015 133.145 ;
        RECT 74.680 133.105 74.880 133.275 ;
        RECT 73.770 133.020 74.170 133.105 ;
        RECT 72.905 132.625 73.165 132.895 ;
        RECT 73.500 132.365 73.670 132.880 ;
        RECT 73.840 132.585 74.170 133.020 ;
        RECT 74.340 132.365 74.510 132.975 ;
        RECT 74.680 132.580 75.010 133.105 ;
        RECT 75.275 132.365 75.485 132.895 ;
        RECT 75.760 132.815 75.930 133.275 ;
        RECT 76.100 133.315 76.420 134.275 ;
        RECT 76.590 133.525 76.780 134.245 ;
        RECT 76.950 133.345 77.120 134.415 ;
        RECT 77.290 134.115 77.460 134.915 ;
        RECT 77.630 134.470 78.735 134.640 ;
        RECT 77.630 133.855 77.800 134.470 ;
        RECT 78.945 134.320 79.195 134.745 ;
        RECT 79.365 134.455 79.630 134.915 ;
        RECT 77.970 133.935 78.500 134.300 ;
        RECT 78.945 134.190 79.250 134.320 ;
        RECT 77.290 133.765 77.800 133.855 ;
        RECT 77.290 133.595 78.160 133.765 ;
        RECT 77.290 133.525 77.460 133.595 ;
        RECT 77.580 133.345 77.780 133.375 ;
        RECT 76.100 132.985 76.565 133.315 ;
        RECT 76.950 133.045 77.780 133.345 ;
        RECT 76.950 132.815 77.120 133.045 ;
        RECT 75.760 132.645 76.545 132.815 ;
        RECT 76.715 132.645 77.120 132.815 ;
        RECT 77.300 132.365 77.670 132.865 ;
        RECT 77.990 132.815 78.160 133.595 ;
        RECT 78.330 133.235 78.500 133.935 ;
        RECT 78.670 133.405 78.910 134.000 ;
        RECT 78.330 133.015 78.855 133.235 ;
        RECT 79.080 133.085 79.250 134.190 ;
        RECT 79.025 132.955 79.250 133.085 ;
        RECT 79.420 132.995 79.700 133.945 ;
        RECT 79.025 132.815 79.195 132.955 ;
        RECT 77.990 132.645 78.665 132.815 ;
        RECT 78.860 132.645 79.195 132.815 ;
        RECT 79.365 132.365 79.615 132.825 ;
        RECT 79.870 132.625 80.055 134.745 ;
        RECT 80.225 134.415 80.555 134.915 ;
        RECT 80.725 134.245 80.895 134.745 ;
        RECT 80.230 134.075 80.895 134.245 ;
        RECT 81.330 134.680 81.540 135.720 ;
        RECT 88.360 135.340 89.270 136.230 ;
        RECT 89.875 135.665 90.045 136.335 ;
        RECT 91.355 136.255 91.605 136.585 ;
        RECT 92.595 136.565 92.765 136.690 ;
        RECT 91.775 136.335 92.765 136.565 ;
        RECT 90.215 136.085 91.195 136.165 ;
        RECT 91.795 136.085 92.425 136.165 ;
        RECT 90.215 135.835 92.425 136.085 ;
        RECT 89.875 135.455 91.185 135.665 ;
        RECT 88.370 135.140 89.260 135.340 ;
        RECT 89.875 135.310 90.045 135.455 ;
        RECT 91.360 135.140 91.600 135.835 ;
        RECT 92.595 135.665 92.765 136.335 ;
        RECT 91.775 135.630 92.765 135.665 ;
        RECT 93.040 136.530 99.780 136.700 ;
        RECT 93.040 135.630 93.210 136.530 ;
        RECT 93.550 135.660 93.720 135.990 ;
        RECT 93.890 135.960 98.930 136.130 ;
        RECT 91.775 135.455 93.210 135.630 ;
        RECT 93.890 135.520 98.930 135.690 ;
        RECT 99.100 135.660 99.270 135.990 ;
        RECT 92.590 135.430 93.210 135.455 ;
        RECT 92.595 135.310 92.765 135.430 ;
        RECT 88.370 134.710 91.610 135.140 ;
        RECT 93.040 135.120 93.210 135.430 ;
        RECT 99.610 135.120 99.780 136.530 ;
        RECT 93.040 134.950 99.780 135.120 ;
        RECT 100.140 135.110 100.310 137.310 ;
        RECT 100.940 136.800 102.940 136.970 ;
        RECT 103.570 136.640 104.490 137.310 ;
        RECT 103.050 136.630 104.490 136.640 ;
        RECT 100.710 135.790 100.880 136.630 ;
        RECT 103.000 135.850 104.490 136.630 ;
        RECT 103.000 135.790 103.170 135.850 ;
        RECT 103.570 135.620 104.490 135.850 ;
        RECT 100.940 135.450 102.940 135.620 ;
        RECT 103.570 135.110 103.740 135.620 ;
        RECT 100.140 134.940 103.740 135.110 ;
        RECT 81.330 134.610 84.000 134.680 ;
        RECT 80.230 133.085 80.460 134.075 ;
        RECT 80.630 133.255 80.980 133.905 ;
        RECT 80.230 132.915 80.895 133.085 ;
        RECT 80.225 132.365 80.555 132.745 ;
        RECT 80.725 132.625 80.895 132.915 ;
        RECT 70.930 132.360 81.070 132.365 ;
        RECT 81.330 132.360 84.500 134.610 ;
        RECT 70.930 132.195 84.500 132.360 ;
        RECT 70.930 132.190 71.520 132.195 ;
        RECT 80.360 132.190 84.500 132.195 ;
        RECT 81.300 131.730 84.500 132.190 ;
        RECT 89.270 131.840 110.850 132.490 ;
        RECT 111.480 131.840 112.920 131.860 ;
        RECT 70.860 131.575 71.640 131.590 ;
        RECT 70.860 131.500 81.130 131.575 ;
        RECT 70.015 131.420 81.130 131.500 ;
        RECT 70.015 131.330 71.250 131.420 ;
        RECT 71.470 131.405 81.130 131.420 ;
        RECT 70.015 130.540 70.185 131.330 ;
        RECT 70.015 130.370 70.860 130.540 ;
        RECT 71.565 130.265 71.815 131.405 ;
        RECT 71.985 130.265 72.320 131.235 ;
        RECT 72.490 130.265 72.705 131.405 ;
        RECT 72.895 130.485 73.225 131.215 ;
        RECT 73.565 130.490 73.740 131.405 ;
        RECT 70.930 128.880 71.260 129.770 ;
        RECT 71.565 128.880 71.815 129.675 ;
        RECT 71.985 129.655 72.200 130.265 ;
        RECT 72.895 130.095 73.165 130.485 ;
        RECT 73.910 130.345 74.240 131.190 ;
        RECT 74.410 130.395 74.580 131.405 ;
        RECT 74.750 130.675 75.090 131.235 ;
        RECT 75.325 130.905 75.640 131.405 ;
        RECT 75.820 130.935 76.705 131.105 ;
        RECT 72.370 129.765 73.165 130.095 ;
        RECT 71.985 129.035 72.240 129.655 ;
        RECT 70.930 128.855 71.815 128.880 ;
        RECT 72.410 128.855 72.740 129.595 ;
        RECT 72.965 129.385 73.165 129.765 ;
        RECT 73.830 130.265 74.240 130.345 ;
        RECT 74.750 130.300 75.650 130.675 ;
        RECT 73.830 130.215 74.065 130.265 ;
        RECT 73.830 129.635 74.020 130.215 ;
        RECT 74.750 130.095 74.940 130.300 ;
        RECT 75.820 130.095 75.990 130.935 ;
        RECT 76.930 130.905 77.180 131.235 ;
        RECT 74.190 129.765 74.940 130.095 ;
        RECT 75.110 129.765 75.990 130.095 ;
        RECT 73.830 129.595 74.075 129.635 ;
        RECT 74.740 129.595 74.940 129.765 ;
        RECT 73.830 129.510 74.230 129.595 ;
        RECT 72.965 129.115 73.225 129.385 ;
        RECT 73.560 128.855 73.730 129.370 ;
        RECT 73.900 129.075 74.230 129.510 ;
        RECT 74.400 128.855 74.570 129.465 ;
        RECT 74.740 129.070 75.070 129.595 ;
        RECT 75.335 128.855 75.545 129.385 ;
        RECT 75.820 129.305 75.990 129.765 ;
        RECT 76.160 129.805 76.480 130.765 ;
        RECT 76.650 130.015 76.840 130.735 ;
        RECT 77.010 129.835 77.180 130.905 ;
        RECT 77.350 130.605 77.520 131.405 ;
        RECT 77.690 130.960 78.795 131.130 ;
        RECT 77.690 130.345 77.860 130.960 ;
        RECT 79.005 130.810 79.255 131.235 ;
        RECT 79.425 130.945 79.690 131.405 ;
        RECT 78.030 130.425 78.560 130.790 ;
        RECT 79.005 130.680 79.310 130.810 ;
        RECT 77.350 130.255 77.860 130.345 ;
        RECT 77.350 130.085 78.220 130.255 ;
        RECT 77.350 130.015 77.520 130.085 ;
        RECT 77.640 129.835 77.840 129.865 ;
        RECT 76.160 129.475 76.625 129.805 ;
        RECT 77.010 129.535 77.840 129.835 ;
        RECT 77.010 129.305 77.180 129.535 ;
        RECT 75.820 129.135 76.605 129.305 ;
        RECT 76.775 129.135 77.180 129.305 ;
        RECT 77.360 128.855 77.730 129.355 ;
        RECT 78.050 129.305 78.220 130.085 ;
        RECT 78.390 129.725 78.560 130.425 ;
        RECT 78.730 129.895 78.970 130.490 ;
        RECT 78.390 129.505 78.915 129.725 ;
        RECT 79.140 129.575 79.310 130.680 ;
        RECT 79.085 129.445 79.310 129.575 ;
        RECT 79.480 129.485 79.760 130.435 ;
        RECT 79.085 129.305 79.255 129.445 ;
        RECT 78.050 129.135 78.725 129.305 ;
        RECT 78.920 129.135 79.255 129.305 ;
        RECT 79.425 128.855 79.675 129.315 ;
        RECT 79.930 129.115 80.115 131.235 ;
        RECT 80.285 130.905 80.615 131.405 ;
        RECT 80.785 130.735 80.955 131.235 ;
        RECT 80.290 130.565 80.955 130.735 ;
        RECT 80.290 129.575 80.520 130.565 ;
        RECT 80.690 129.745 81.040 130.395 ;
        RECT 80.290 129.405 80.955 129.575 ;
        RECT 80.285 128.860 80.615 129.235 ;
        RECT 80.785 129.115 80.955 129.405 ;
        RECT 81.300 128.860 83.560 131.730 ;
        RECT 84.750 131.670 112.920 131.840 ;
        RECT 84.750 129.300 84.920 131.670 ;
        RECT 85.400 129.780 87.560 131.190 ;
        RECT 108.820 129.780 110.980 131.190 ;
        RECT 111.460 129.300 112.920 131.670 ;
        RECT 84.750 129.160 112.920 129.300 ;
        RECT 84.750 129.130 111.630 129.160 ;
        RECT 80.285 128.855 83.560 128.860 ;
        RECT 70.930 128.720 83.560 128.855 ;
        RECT 70.930 128.690 82.630 128.720 ;
        RECT 71.470 128.685 82.630 128.690 ;
        RECT 80.410 128.680 82.630 128.685 ;
        RECT 81.300 128.670 81.550 128.680 ;
        RECT 82.420 128.670 82.630 128.680 ;
        RECT 151.870 29.320 152.970 29.530 ;
        RECT 106.250 28.260 109.740 28.430 ;
        RECT 106.250 27.510 106.420 28.260 ;
        RECT 107.050 27.750 107.850 27.920 ;
        RECT 108.140 27.750 108.940 27.920 ;
        RECT 106.220 26.860 106.510 27.510 ;
        RECT 106.250 23.520 106.420 26.860 ;
        RECT 106.820 24.245 106.990 27.535 ;
        RECT 107.910 24.245 108.080 27.535 ;
        RECT 109.000 24.245 109.170 27.535 ;
        RECT 107.050 23.860 107.850 24.030 ;
        RECT 108.140 23.860 108.940 24.030 ;
        RECT 109.570 23.520 109.740 28.260 ;
        RECT 111.370 28.260 114.860 28.430 ;
        RECT 111.370 27.400 111.540 28.260 ;
        RECT 112.170 27.750 112.970 27.920 ;
        RECT 113.260 27.750 114.060 27.920 ;
        RECT 111.320 26.700 111.610 27.400 ;
        RECT 106.250 23.350 109.740 23.520 ;
        RECT 111.370 23.520 111.540 26.700 ;
        RECT 111.940 24.245 112.110 27.535 ;
        RECT 113.030 24.245 113.200 27.535 ;
        RECT 114.120 24.245 114.290 27.535 ;
        RECT 112.170 23.860 112.970 24.030 ;
        RECT 113.260 23.860 114.060 24.030 ;
        RECT 114.690 23.520 114.860 28.260 ;
        RECT 116.490 28.250 119.980 28.420 ;
        RECT 116.490 27.390 116.660 28.250 ;
        RECT 117.290 27.740 118.090 27.910 ;
        RECT 118.380 27.740 119.180 27.910 ;
        RECT 116.480 26.770 116.670 27.390 ;
        RECT 111.370 23.350 114.860 23.520 ;
        RECT 116.490 23.510 116.660 26.770 ;
        RECT 117.060 24.235 117.230 27.525 ;
        RECT 118.150 24.235 118.320 27.525 ;
        RECT 119.240 24.235 119.410 27.525 ;
        RECT 117.290 23.850 118.090 24.020 ;
        RECT 118.380 23.850 119.180 24.020 ;
        RECT 119.810 23.510 119.980 28.250 ;
        RECT 121.610 28.250 125.100 28.420 ;
        RECT 121.610 27.470 121.780 28.250 ;
        RECT 122.410 27.740 123.210 27.910 ;
        RECT 123.500 27.740 124.300 27.910 ;
        RECT 121.570 26.820 121.800 27.470 ;
        RECT 116.490 23.340 119.980 23.510 ;
        RECT 121.610 23.510 121.780 26.820 ;
        RECT 122.180 24.235 122.350 27.525 ;
        RECT 123.270 24.235 123.440 27.525 ;
        RECT 124.360 24.235 124.530 27.525 ;
        RECT 122.410 23.850 123.210 24.020 ;
        RECT 123.500 23.850 124.300 24.020 ;
        RECT 124.930 23.510 125.100 28.250 ;
        RECT 143.230 27.820 145.210 28.410 ;
        RECT 151.870 28.090 153.640 29.320 ;
        RECT 152.970 27.820 153.640 28.090 ;
        RECT 121.610 23.340 125.100 23.510 ;
        RECT 139.030 27.580 142.110 27.590 ;
        RECT 143.700 27.580 144.950 27.820 ;
        RECT 139.030 27.420 144.950 27.580 ;
        RECT 121.570 22.190 125.060 22.360 ;
        RECT 99.400 21.610 102.150 21.780 ;
        RECT 99.400 20.860 99.570 21.610 ;
        RECT 100.610 21.100 100.940 21.270 ;
        RECT 99.300 20.430 99.620 20.860 ;
        RECT 99.400 18.120 99.570 20.430 ;
        RECT 99.970 18.845 100.140 20.885 ;
        RECT 100.450 18.845 100.620 20.885 ;
        RECT 100.930 18.845 101.100 20.885 ;
        RECT 101.410 18.845 101.580 20.885 ;
        RECT 100.130 18.460 100.460 18.630 ;
        RECT 101.090 18.460 101.420 18.630 ;
        RECT 101.980 18.120 102.150 21.610 ;
        RECT 103.790 21.550 108.220 21.720 ;
        RECT 103.790 20.830 103.960 21.550 ;
        RECT 104.590 21.040 105.340 21.210 ;
        RECT 105.630 21.040 106.380 21.210 ;
        RECT 106.670 21.040 107.420 21.210 ;
        RECT 103.780 20.400 103.980 20.830 ;
        RECT 99.400 17.950 102.150 18.120 ;
        RECT 103.790 18.060 103.960 20.400 ;
        RECT 104.360 18.785 104.530 20.825 ;
        RECT 105.400 18.785 105.570 20.825 ;
        RECT 106.440 18.785 106.610 20.825 ;
        RECT 107.480 18.785 107.650 20.825 ;
        RECT 104.590 18.400 105.340 18.570 ;
        RECT 105.630 18.400 106.380 18.570 ;
        RECT 106.670 18.400 107.420 18.570 ;
        RECT 108.050 18.060 108.220 21.550 ;
        RECT 109.850 21.550 114.280 21.720 ;
        RECT 109.850 20.790 110.020 21.550 ;
        RECT 110.650 21.040 111.400 21.210 ;
        RECT 111.690 21.040 112.440 21.210 ;
        RECT 112.730 21.040 113.480 21.210 ;
        RECT 109.810 20.380 110.080 20.790 ;
        RECT 103.790 17.890 108.220 18.060 ;
        RECT 109.850 18.060 110.020 20.380 ;
        RECT 110.420 18.785 110.590 20.825 ;
        RECT 111.460 18.785 111.630 20.825 ;
        RECT 112.500 18.785 112.670 20.825 ;
        RECT 113.540 18.785 113.710 20.825 ;
        RECT 110.650 18.400 111.400 18.570 ;
        RECT 111.690 18.400 112.440 18.570 ;
        RECT 112.730 18.400 113.480 18.570 ;
        RECT 114.110 18.060 114.280 21.550 ;
        RECT 115.910 21.540 120.340 21.710 ;
        RECT 115.910 20.770 116.080 21.540 ;
        RECT 116.710 21.030 117.460 21.200 ;
        RECT 117.750 21.030 118.500 21.200 ;
        RECT 118.790 21.030 119.540 21.200 ;
        RECT 115.850 20.230 116.110 20.770 ;
        RECT 109.850 17.890 114.280 18.060 ;
        RECT 115.910 18.050 116.080 20.230 ;
        RECT 116.480 18.775 116.650 20.815 ;
        RECT 117.520 18.775 117.690 20.815 ;
        RECT 118.560 18.775 118.730 20.815 ;
        RECT 119.600 18.775 119.770 20.815 ;
        RECT 116.710 18.390 117.460 18.560 ;
        RECT 117.750 18.390 118.500 18.560 ;
        RECT 118.790 18.390 119.540 18.560 ;
        RECT 120.170 18.050 120.340 21.540 ;
        RECT 121.570 19.090 121.740 22.190 ;
        RECT 122.370 21.680 123.170 21.850 ;
        RECT 123.460 21.680 124.260 21.850 ;
        RECT 121.510 18.320 121.790 19.090 ;
        RECT 115.910 17.880 120.340 18.050 ;
        RECT 121.570 17.540 121.740 18.320 ;
        RECT 122.140 18.220 122.310 21.510 ;
        RECT 123.230 18.220 123.400 21.510 ;
        RECT 124.320 18.220 124.490 21.510 ;
        RECT 122.370 17.880 123.170 18.050 ;
        RECT 123.460 17.880 124.260 18.050 ;
        RECT 124.890 17.540 125.060 22.190 ;
        RECT 139.030 19.930 139.200 27.420 ;
        RECT 141.830 27.270 144.950 27.420 ;
        RECT 151.060 27.650 153.640 27.820 ;
        RECT 141.830 27.100 146.680 27.270 ;
        RECT 139.815 26.910 140.145 27.080 ;
        RECT 140.405 26.910 140.735 27.080 ;
        RECT 140.995 26.910 141.325 27.080 ;
        RECT 141.830 26.790 144.950 27.100 ;
        RECT 139.600 20.655 139.770 26.695 ;
        RECT 140.190 20.655 140.360 26.695 ;
        RECT 140.780 20.655 140.950 26.695 ;
        RECT 141.370 20.655 141.540 26.695 ;
        RECT 141.830 26.220 144.970 26.790 ;
        RECT 145.565 26.590 145.895 26.760 ;
        RECT 139.815 20.270 140.145 20.440 ;
        RECT 140.405 20.270 140.735 20.440 ;
        RECT 140.995 20.270 141.325 20.440 ;
        RECT 141.940 19.930 142.110 26.220 ;
        RECT 143.710 26.180 144.970 26.220 ;
        RECT 139.030 19.760 142.110 19.930 ;
        RECT 144.780 19.610 144.950 26.180 ;
        RECT 145.350 20.335 145.520 26.375 ;
        RECT 145.940 20.335 146.110 26.375 ;
        RECT 145.565 19.950 145.895 20.120 ;
        RECT 146.510 19.610 146.680 27.100 ;
        RECT 144.780 19.440 146.680 19.610 ;
        RECT 151.060 19.160 151.230 27.650 ;
        RECT 151.845 27.140 152.175 27.310 ;
        RECT 152.435 27.140 152.765 27.310 ;
        RECT 152.970 27.170 153.640 27.650 ;
        RECT 151.630 19.885 151.800 26.925 ;
        RECT 152.220 19.885 152.390 26.925 ;
        RECT 152.810 19.885 152.980 26.925 ;
        RECT 151.845 19.500 152.175 19.670 ;
        RECT 152.435 19.500 152.765 19.670 ;
        RECT 153.380 19.160 153.550 27.170 ;
        RECT 151.060 18.990 153.550 19.160 ;
        RECT 140.995 18.225 142.895 18.395 ;
        RECT 121.570 17.370 125.060 17.540 ;
        RECT 137.245 17.765 139.145 17.935 ;
        RECT 99.770 16.820 102.040 16.990 ;
        RECT 99.770 14.440 99.940 16.820 ;
        RECT 100.500 16.310 100.830 16.480 ;
        RECT 99.730 13.920 100.000 14.440 ;
        RECT 99.770 13.170 99.940 13.920 ;
        RECT 100.340 13.850 100.510 16.140 ;
        RECT 100.820 13.850 100.990 16.140 ;
        RECT 101.300 13.850 101.470 16.140 ;
        RECT 100.980 13.510 101.310 13.680 ;
        RECT 101.870 13.170 102.040 16.820 ;
        RECT 104.570 16.890 107.960 17.060 ;
        RECT 104.570 14.600 104.740 16.890 ;
        RECT 105.370 16.380 106.120 16.550 ;
        RECT 106.410 16.380 107.160 16.550 ;
        RECT 104.550 14.010 104.740 14.600 ;
        RECT 99.770 13.000 102.040 13.170 ;
        RECT 104.570 13.240 104.740 14.010 ;
        RECT 105.140 13.920 105.310 16.210 ;
        RECT 106.180 13.920 106.350 16.210 ;
        RECT 107.220 13.920 107.390 16.210 ;
        RECT 105.370 13.580 106.120 13.750 ;
        RECT 106.410 13.580 107.160 13.750 ;
        RECT 107.790 13.240 107.960 16.890 ;
        RECT 104.570 13.070 107.960 13.240 ;
        RECT 110.660 16.870 114.050 17.040 ;
        RECT 110.660 14.530 110.830 16.870 ;
        RECT 111.460 16.360 112.210 16.530 ;
        RECT 112.500 16.360 113.250 16.530 ;
        RECT 110.660 13.970 110.840 14.530 ;
        RECT 110.660 13.220 110.830 13.970 ;
        RECT 111.230 13.900 111.400 16.190 ;
        RECT 112.270 13.900 112.440 16.190 ;
        RECT 113.310 13.900 113.480 16.190 ;
        RECT 111.460 13.560 112.210 13.730 ;
        RECT 112.500 13.560 113.250 13.730 ;
        RECT 113.880 13.220 114.050 16.870 ;
        RECT 116.670 16.880 120.060 17.050 ;
        RECT 116.670 14.470 116.840 16.880 ;
        RECT 117.470 16.370 118.220 16.540 ;
        RECT 118.510 16.370 119.260 16.540 ;
        RECT 116.600 13.970 116.870 14.470 ;
        RECT 110.660 13.050 114.050 13.220 ;
        RECT 116.670 13.230 116.840 13.970 ;
        RECT 117.240 13.910 117.410 16.200 ;
        RECT 118.280 13.910 118.450 16.200 ;
        RECT 119.320 13.910 119.490 16.200 ;
        RECT 117.470 13.570 118.220 13.740 ;
        RECT 118.510 13.570 119.260 13.740 ;
        RECT 119.890 13.230 120.060 16.880 ;
        RECT 137.245 14.365 137.415 17.765 ;
        RECT 138.030 17.255 138.360 17.425 ;
        RECT 137.815 15.045 137.985 17.085 ;
        RECT 138.405 15.045 138.575 17.085 ;
        RECT 138.030 14.705 138.360 14.875 ;
        RECT 138.975 14.365 139.145 17.765 ;
        RECT 140.995 14.840 141.165 18.225 ;
        RECT 141.780 17.715 142.110 17.885 ;
        RECT 141.565 15.505 141.735 17.545 ;
        RECT 142.155 15.505 142.325 17.545 ;
        RECT 141.780 15.165 142.110 15.335 ;
        RECT 140.940 14.825 141.720 14.840 ;
        RECT 142.725 14.825 142.895 18.225 ;
        RECT 151.080 17.350 152.130 18.990 ;
        RECT 150.465 17.180 154.065 17.350 ;
        RECT 140.940 14.655 142.895 14.825 ;
        RECT 144.280 16.260 146.380 16.430 ;
        RECT 140.940 14.400 141.670 14.655 ;
        RECT 137.245 14.360 139.145 14.365 ;
        RECT 137.220 14.195 139.145 14.360 ;
        RECT 140.930 14.340 141.670 14.400 ;
        RECT 141.910 14.340 142.370 14.380 ;
        RECT 137.220 13.980 137.840 14.195 ;
        RECT 140.930 14.070 142.370 14.340 ;
        RECT 144.280 14.200 144.450 16.260 ;
        RECT 145.080 15.750 145.580 15.920 ;
        RECT 144.850 14.840 145.020 15.580 ;
        RECT 145.640 14.840 145.810 15.580 ;
        RECT 145.080 14.500 145.580 14.670 ;
        RECT 144.280 14.160 144.870 14.200 ;
        RECT 146.210 14.160 146.380 16.260 ;
        RECT 150.465 14.690 150.635 17.180 ;
        RECT 151.265 16.670 153.265 16.840 ;
        RECT 151.035 15.415 151.205 16.455 ;
        RECT 153.325 15.415 153.495 16.455 ;
        RECT 151.265 15.030 153.265 15.200 ;
        RECT 153.895 14.690 154.065 17.180 ;
        RECT 150.465 14.520 154.065 14.690 ;
        RECT 137.220 13.820 138.020 13.980 ;
        RECT 140.930 13.970 142.210 14.070 ;
        RECT 144.280 13.990 146.380 14.160 ;
        RECT 140.930 13.960 141.520 13.970 ;
        RECT 137.220 13.640 138.630 13.820 ;
        RECT 144.300 13.740 144.870 13.990 ;
        RECT 116.670 13.060 120.060 13.230 ;
        RECT 137.190 13.200 138.630 13.640 ;
        RECT 138.000 13.100 138.630 13.200 ;
        RECT 143.990 13.180 145.070 13.740 ;
        RECT 148.760 13.290 155.360 13.370 ;
        RECT 145.830 13.200 155.360 13.290 ;
        RECT 145.830 12.770 148.960 13.200 ;
        RECT 146.030 12.690 148.960 12.770 ;
        RECT 149.560 12.690 154.560 12.860 ;
        RECT 104.530 12.030 108.020 12.200 ;
        RECT 104.530 8.950 104.700 12.030 ;
        RECT 105.330 11.520 106.130 11.690 ;
        RECT 106.420 11.520 107.220 11.690 ;
        RECT 104.480 8.110 104.780 8.950 ;
        RECT 104.530 7.380 104.700 8.110 ;
        RECT 105.100 8.060 105.270 11.350 ;
        RECT 106.190 8.060 106.360 11.350 ;
        RECT 107.280 8.060 107.450 11.350 ;
        RECT 105.330 7.720 106.130 7.890 ;
        RECT 106.420 7.720 107.220 7.890 ;
        RECT 107.850 7.380 108.020 12.030 ;
        RECT 110.630 12.030 114.120 12.200 ;
        RECT 110.630 8.970 110.800 12.030 ;
        RECT 111.430 11.520 112.230 11.690 ;
        RECT 112.520 11.520 113.320 11.690 ;
        RECT 110.510 8.130 110.810 8.970 ;
        RECT 104.530 7.210 108.020 7.380 ;
        RECT 110.630 7.380 110.800 8.130 ;
        RECT 111.200 8.060 111.370 11.350 ;
        RECT 112.290 8.060 112.460 11.350 ;
        RECT 113.380 8.060 113.550 11.350 ;
        RECT 111.430 7.720 112.230 7.890 ;
        RECT 112.520 7.720 113.320 7.890 ;
        RECT 113.950 7.380 114.120 12.030 ;
        RECT 116.710 12.050 120.200 12.220 ;
        RECT 116.710 8.820 116.880 12.050 ;
        RECT 117.510 11.540 118.310 11.710 ;
        RECT 118.600 11.540 119.400 11.710 ;
        RECT 116.660 8.170 116.930 8.820 ;
        RECT 110.630 7.210 114.120 7.380 ;
        RECT 116.710 7.400 116.880 8.170 ;
        RECT 117.280 8.080 117.450 11.370 ;
        RECT 118.370 8.080 118.540 11.370 ;
        RECT 119.460 8.080 119.630 11.370 ;
        RECT 117.510 7.740 118.310 7.910 ;
        RECT 118.600 7.740 119.400 7.910 ;
        RECT 120.030 7.400 120.200 12.050 ;
        RECT 148.760 10.800 148.930 12.690 ;
        RECT 149.330 11.480 149.500 12.520 ;
        RECT 154.620 11.480 154.790 12.520 ;
        RECT 149.560 11.140 154.560 11.310 ;
        RECT 155.190 10.800 155.360 13.200 ;
        RECT 148.760 10.630 155.360 10.800 ;
        RECT 116.710 7.230 120.200 7.400 ;
      LAYER met1 ;
        RECT 42.070 223.290 43.670 224.310 ;
        RECT 45.430 223.360 48.390 223.680 ;
        RECT 7.700 222.130 8.860 222.150 ;
        RECT 6.740 221.310 9.860 222.130 ;
        RECT 7.700 213.140 8.860 221.310 ;
        RECT 43.110 221.070 43.410 223.290 ;
        RECT 45.480 221.070 45.780 223.360 ;
        RECT 51.920 221.070 63.400 221.360 ;
        RECT 54.490 221.060 63.400 221.070 ;
        RECT 60.740 221.040 63.400 221.060 ;
        RECT 60.750 220.890 63.300 221.040 ;
        RECT 17.200 214.780 17.760 214.810 ;
        RECT 18.190 214.780 18.690 214.850 ;
        RECT 17.200 214.540 18.690 214.780 ;
        RECT 30.900 214.720 31.670 215.430 ;
        RECT 17.200 214.500 17.760 214.540 ;
        RECT 18.190 214.440 18.690 214.540 ;
        RECT 30.030 214.340 31.670 214.720 ;
        RECT 41.910 214.800 42.970 214.810 ;
        RECT 43.110 214.800 43.410 220.770 ;
        RECT 45.480 216.490 45.780 220.770 ;
        RECT 44.340 215.950 45.840 216.490 ;
        RECT 41.910 214.460 43.410 214.800 ;
        RECT 46.860 214.750 47.430 217.620 ;
        RECT 42.850 214.390 43.410 214.460 ;
        RECT 42.850 214.380 43.400 214.390 ;
        RECT 30.540 214.330 31.670 214.340 ;
        RECT 23.220 214.180 31.960 214.190 ;
        RECT 35.130 214.180 43.870 214.190 ;
        RECT 10.420 214.060 43.870 214.180 ;
        RECT 44.070 214.060 46.460 214.160 ;
        RECT 10.420 213.830 46.460 214.060 ;
        RECT 10.420 213.720 43.870 213.830 ;
        RECT 10.420 213.700 19.160 213.720 ;
        RECT 17.300 213.530 17.600 213.540 ;
        RECT 17.270 213.160 17.690 213.530 ;
        RECT 19.460 213.490 19.760 213.720 ;
        RECT 23.220 213.710 31.960 213.720 ;
        RECT 30.090 213.550 30.420 213.560 ;
        RECT 19.450 213.210 19.770 213.490 ;
        RECT 30.060 213.170 30.510 213.550 ;
        RECT 32.200 213.310 32.620 213.720 ;
        RECT 35.130 213.710 43.870 213.720 ;
        RECT 41.990 213.560 42.320 213.570 ;
        RECT 32.260 213.150 32.580 213.310 ;
        RECT 41.970 213.230 42.410 213.560 ;
        RECT 7.620 212.910 8.890 213.140 ;
        RECT 18.860 212.910 19.030 212.920 ;
        RECT 7.620 212.580 10.850 212.910 ;
        RECT 11.800 212.880 12.160 212.900 ;
        RECT 11.790 212.870 12.160 212.880 ;
        RECT 18.540 212.870 19.030 212.910 ;
        RECT 11.790 212.840 19.030 212.870 ;
        RECT 23.310 212.840 23.630 212.940 ;
        RECT 24.590 212.930 24.970 212.970 ;
        RECT 11.790 212.690 23.630 212.840 ;
        RECT 11.790 212.630 12.160 212.690 ;
        RECT 18.540 212.640 23.630 212.690 ;
        RECT 24.570 212.920 24.970 212.930 ;
        RECT 30.890 212.920 31.870 212.970 ;
        RECT 36.500 212.950 36.950 212.990 ;
        RECT 42.810 212.960 43.230 213.030 ;
        RECT 42.810 212.950 43.750 212.960 ;
        RECT 24.570 212.890 31.870 212.920 ;
        RECT 35.150 212.890 35.550 212.920 ;
        RECT 24.570 212.690 35.550 212.890 ;
        RECT 24.570 212.650 24.970 212.690 ;
        RECT 11.800 212.620 12.160 212.630 ;
        RECT 7.620 211.980 8.890 212.580 ;
        RECT 11.385 212.480 11.675 212.525 ;
        RECT 12.575 212.480 12.865 212.525 ;
        RECT 15.095 212.480 15.385 212.525 ;
        RECT 18.860 212.480 19.030 212.640 ;
        RECT 23.310 212.540 23.630 212.640 ;
        RECT 24.590 212.630 24.970 212.650 ;
        RECT 30.890 212.620 35.550 212.690 ;
        RECT 36.500 212.730 43.750 212.950 ;
        RECT 36.500 212.640 36.950 212.730 ;
        RECT 42.810 212.710 43.750 212.730 ;
        RECT 44.070 212.720 46.460 213.830 ;
        RECT 42.810 212.660 43.230 212.710 ;
        RECT 31.620 212.560 35.550 212.620 ;
        RECT 24.185 212.490 24.475 212.535 ;
        RECT 25.375 212.490 25.665 212.535 ;
        RECT 27.895 212.490 28.185 212.535 ;
        RECT 11.385 212.340 15.385 212.480 ;
        RECT 11.385 212.295 11.675 212.340 ;
        RECT 12.575 212.295 12.865 212.340 ;
        RECT 15.095 212.295 15.385 212.340 ;
        RECT 18.760 212.200 19.110 212.480 ;
        RECT 24.185 212.350 28.185 212.490 ;
        RECT 31.620 212.460 31.900 212.560 ;
        RECT 24.185 212.305 24.475 212.350 ;
        RECT 25.375 212.305 25.665 212.350 ;
        RECT 27.895 212.305 28.185 212.350 ;
        RECT 31.570 212.400 31.900 212.460 ;
        RECT 36.095 212.490 36.385 212.535 ;
        RECT 37.285 212.490 37.575 212.535 ;
        RECT 39.805 212.490 40.095 212.535 ;
        RECT 31.570 212.210 31.890 212.400 ;
        RECT 36.095 212.350 40.095 212.490 ;
        RECT 43.530 212.460 43.750 212.710 ;
        RECT 36.095 212.305 36.385 212.350 ;
        RECT 37.285 212.305 37.575 212.350 ;
        RECT 39.805 212.305 40.095 212.350 ;
        RECT 43.490 212.220 43.800 212.460 ;
        RECT 10.990 212.140 11.280 212.185 ;
        RECT 13.090 212.140 13.380 212.185 ;
        RECT 14.660 212.140 14.950 212.185 ;
        RECT 10.990 212.000 14.950 212.140 ;
        RECT 18.860 212.110 19.030 212.200 ;
        RECT 23.790 212.150 24.080 212.195 ;
        RECT 25.890 212.150 26.180 212.195 ;
        RECT 27.460 212.150 27.750 212.195 ;
        RECT 31.620 212.190 31.860 212.210 ;
        RECT 10.990 211.955 11.280 212.000 ;
        RECT 13.090 211.955 13.380 212.000 ;
        RECT 14.660 211.955 14.950 212.000 ;
        RECT 23.790 212.010 27.750 212.150 ;
        RECT 23.790 211.965 24.080 212.010 ;
        RECT 25.890 211.965 26.180 212.010 ;
        RECT 27.460 211.965 27.750 212.010 ;
        RECT 35.700 212.150 35.990 212.195 ;
        RECT 37.800 212.150 38.090 212.195 ;
        RECT 39.370 212.150 39.660 212.195 ;
        RECT 35.700 212.010 39.660 212.150 ;
        RECT 43.530 212.110 43.750 212.220 ;
        RECT 35.700 211.965 35.990 212.010 ;
        RECT 37.800 211.965 38.090 212.010 ;
        RECT 39.370 211.965 39.660 212.010 ;
        RECT 9.120 211.010 43.870 211.470 ;
        RECT 9.140 210.980 19.160 211.010 ;
        RECT 23.220 210.990 31.960 211.010 ;
        RECT 35.130 210.990 43.870 211.010 ;
        RECT 9.140 209.060 11.990 210.980 ;
        RECT 9.070 206.560 12.260 209.060 ;
        RECT 21.960 208.790 22.960 208.820 ;
        RECT 19.220 206.880 25.350 208.790 ;
        RECT 18.150 202.820 19.150 203.820 ;
        RECT 21.960 203.540 22.960 206.880 ;
        RECT 46.960 205.790 47.260 214.750 ;
        RECT 30.960 205.490 47.260 205.790 ;
        RECT 30.960 203.790 31.260 205.490 ;
        RECT 52.220 203.830 52.760 220.770 ;
        RECT 77.370 220.750 78.370 221.750 ;
        RECT 57.410 220.280 78.370 220.750 ;
        RECT 136.590 220.740 137.590 220.760 ;
        RECT 57.410 220.270 65.420 220.280 ;
        RECT 65.800 220.270 78.370 220.280 ;
        RECT 54.960 219.340 56.190 220.260 ;
        RECT 70.585 219.730 70.875 219.775 ;
        RECT 73.705 219.730 73.995 219.775 ;
        RECT 75.595 219.730 75.885 219.775 ;
        RECT 70.585 219.590 75.885 219.730 ;
        RECT 70.585 219.545 70.875 219.590 ;
        RECT 73.705 219.545 73.995 219.590 ;
        RECT 75.595 219.545 75.885 219.590 ;
        RECT 54.960 218.740 57.930 219.340 ;
        RECT 65.000 218.820 65.360 219.150 ;
        RECT 67.360 219.120 67.660 219.170 ;
        RECT 67.290 218.810 67.730 219.120 ;
        RECT 69.280 219.070 69.710 219.180 ;
        RECT 69.280 218.900 69.795 219.070 ;
        RECT 67.360 218.760 67.660 218.810 ;
        RECT 69.505 218.755 69.795 218.900 ;
        RECT 70.585 219.050 70.875 219.095 ;
        RECT 74.165 219.050 74.455 219.095 ;
        RECT 76.000 219.050 76.290 219.095 ;
        RECT 70.585 218.910 76.290 219.050 ;
        RECT 70.585 218.865 70.875 218.910 ;
        RECT 74.165 218.865 74.455 218.910 ;
        RECT 76.000 218.865 76.290 218.910 ;
        RECT 76.470 218.770 77.200 219.110 ;
        RECT 54.960 218.640 56.190 218.740 ;
        RECT 69.205 218.710 69.795 218.755 ;
        RECT 72.445 218.710 73.095 218.755 ;
        RECT 55.100 218.620 56.100 218.640 ;
        RECT 69.205 218.570 73.095 218.710 ;
        RECT 69.205 218.525 69.495 218.570 ;
        RECT 72.445 218.525 73.095 218.570 ;
        RECT 56.400 217.550 77.300 218.030 ;
        RECT 77.710 217.650 78.370 220.270 ;
        RECT 135.950 219.760 137.590 220.740 ;
        RECT 79.070 219.460 80.070 219.570 ;
        RECT 79.070 218.920 111.250 219.460 ;
        RECT 135.950 219.400 136.320 219.760 ;
        RECT 79.070 218.570 80.070 218.920 ;
        RECT 56.400 214.690 57.060 217.550 ;
        RECT 77.620 217.410 78.430 217.650 ;
        RECT 63.580 216.930 78.430 217.410 ;
        RECT 68.610 215.980 68.920 216.020 ;
        RECT 63.830 215.530 64.270 215.840 ;
        RECT 64.530 215.530 64.970 215.840 ;
        RECT 65.760 215.520 66.830 215.780 ;
        RECT 68.610 215.480 69.290 215.980 ;
        RECT 68.610 215.430 68.920 215.480 ;
        RECT 56.400 214.210 69.020 214.690 ;
        RECT 54.160 212.870 55.660 212.890 ;
        RECT 54.160 212.690 56.100 212.870 ;
        RECT 54.160 212.090 56.150 212.690 ;
        RECT 54.160 211.870 56.100 212.090 ;
        RECT 54.160 211.840 55.660 211.870 ;
        RECT 21.950 203.120 22.960 203.540 ;
        RECT 8.000 201.300 8.910 202.790 ;
        RECT 21.950 202.620 22.950 203.120 ;
        RECT 30.560 202.790 31.560 203.790 ;
        RECT 42.940 203.290 52.760 203.830 ;
        RECT 56.400 211.350 57.060 214.210 ;
        RECT 77.620 214.070 78.430 216.930 ;
        RECT 128.380 217.060 129.300 217.130 ;
        RECT 131.750 217.120 132.750 217.220 ;
        RECT 131.750 217.060 132.920 217.120 ;
        RECT 128.380 216.360 132.920 217.060 ;
        RECT 128.380 216.300 132.750 216.360 ;
        RECT 128.380 216.230 129.300 216.300 ;
        RECT 131.750 216.220 132.750 216.300 ;
        RECT 59.670 213.760 78.430 214.070 ;
        RECT 59.670 213.600 78.370 213.760 ;
        RECT 60.630 213.590 62.930 213.600 ;
        RECT 63.310 213.590 65.610 213.600 ;
        RECT 65.800 213.590 78.370 213.600 ;
        RECT 70.585 213.050 70.875 213.095 ;
        RECT 73.705 213.050 73.995 213.095 ;
        RECT 75.595 213.050 75.885 213.095 ;
        RECT 70.585 212.910 75.885 213.050 ;
        RECT 70.585 212.865 70.875 212.910 ;
        RECT 73.705 212.865 73.995 212.910 ;
        RECT 75.595 212.865 75.885 212.910 ;
        RECT 59.440 212.090 60.820 212.690 ;
        RECT 65.250 212.420 65.480 212.470 ;
        RECT 67.390 212.440 67.620 212.460 ;
        RECT 65.190 212.110 65.550 212.420 ;
        RECT 67.290 212.130 67.730 212.440 ;
        RECT 69.280 212.390 69.710 212.520 ;
        RECT 69.280 212.240 69.795 212.390 ;
        RECT 67.390 212.110 67.620 212.130 ;
        RECT 60.010 212.070 60.820 212.090 ;
        RECT 69.505 212.075 69.795 212.240 ;
        RECT 70.585 212.370 70.875 212.415 ;
        RECT 74.165 212.370 74.455 212.415 ;
        RECT 76.000 212.370 76.290 212.415 ;
        RECT 70.585 212.230 76.290 212.370 ;
        RECT 70.585 212.185 70.875 212.230 ;
        RECT 74.165 212.185 74.455 212.230 ;
        RECT 76.000 212.185 76.290 212.230 ;
        RECT 76.430 212.100 76.880 212.500 ;
        RECT 69.205 212.030 69.795 212.075 ;
        RECT 72.445 212.030 73.095 212.075 ;
        RECT 69.205 211.890 73.095 212.030 ;
        RECT 69.205 211.845 69.495 211.890 ;
        RECT 72.445 211.845 73.095 211.890 ;
        RECT 56.400 210.870 77.300 211.350 ;
        RECT 42.940 202.830 43.940 203.290 ;
        RECT 11.130 202.600 36.020 202.620 ;
        RECT 11.130 202.150 45.540 202.600 ;
        RECT 11.130 202.140 33.220 202.150 ;
        RECT 11.130 202.120 33.190 202.140 ;
        RECT 35.880 202.120 45.540 202.150 ;
        RECT 56.400 202.060 57.400 210.870 ;
        RECT 77.710 209.110 78.370 213.590 ;
        RECT 106.380 213.110 108.070 213.810 ;
        RECT 79.040 212.590 108.070 213.110 ;
        RECT 79.020 212.450 108.070 212.590 ;
        RECT 79.020 211.850 80.070 212.450 ;
        RECT 106.380 212.240 108.070 212.450 ;
        RECT 79.070 211.740 80.070 211.850 ;
        RECT 75.250 206.680 78.440 209.110 ;
        RECT 77.710 206.600 78.370 206.680 ;
        RECT 82.120 206.660 84.040 209.000 ;
        RECT 11.710 201.600 12.000 201.645 ;
        RECT 13.810 201.600 14.100 201.645 ;
        RECT 15.380 201.600 15.670 201.645 ;
        RECT 11.710 201.460 15.670 201.600 ;
        RECT 11.710 201.415 12.000 201.460 ;
        RECT 13.810 201.415 14.100 201.460 ;
        RECT 15.380 201.415 15.670 201.460 ;
        RECT 24.130 201.600 24.420 201.645 ;
        RECT 26.230 201.600 26.520 201.645 ;
        RECT 27.800 201.600 28.090 201.645 ;
        RECT 24.130 201.460 28.090 201.600 ;
        RECT 24.130 201.415 24.420 201.460 ;
        RECT 26.230 201.415 26.520 201.460 ;
        RECT 27.800 201.415 28.090 201.460 ;
        RECT 36.450 201.580 36.740 201.625 ;
        RECT 38.550 201.580 38.840 201.625 ;
        RECT 40.120 201.580 40.410 201.625 ;
        RECT 36.450 201.440 40.410 201.580 ;
        RECT 36.450 201.395 36.740 201.440 ;
        RECT 38.550 201.395 38.840 201.440 ;
        RECT 40.120 201.395 40.410 201.440 ;
        RECT 8.000 201.050 10.770 201.300 ;
        RECT 12.105 201.260 12.395 201.305 ;
        RECT 13.295 201.260 13.585 201.305 ;
        RECT 15.815 201.260 16.105 201.305 ;
        RECT 12.105 201.120 16.105 201.260 ;
        RECT 11.250 201.050 11.560 201.120 ;
        RECT 12.105 201.075 12.395 201.120 ;
        RECT 13.295 201.075 13.585 201.120 ;
        RECT 15.815 201.075 16.105 201.120 ;
        RECT 8.000 200.650 11.560 201.050 ;
        RECT 20.050 200.940 20.280 200.990 ;
        RECT 23.620 200.940 24.010 201.320 ;
        RECT 24.525 201.260 24.815 201.305 ;
        RECT 25.715 201.260 26.005 201.305 ;
        RECT 28.235 201.260 28.525 201.305 ;
        RECT 24.525 201.120 28.525 201.260 ;
        RECT 36.845 201.240 37.135 201.285 ;
        RECT 38.035 201.240 38.325 201.285 ;
        RECT 40.555 201.240 40.845 201.285 ;
        RECT 24.525 201.075 24.815 201.120 ;
        RECT 25.715 201.075 26.005 201.120 ;
        RECT 28.235 201.075 28.525 201.120 ;
        RECT 20.050 200.920 24.010 200.940 ;
        RECT 8.000 200.300 10.770 200.650 ;
        RECT 12.500 200.640 24.010 200.920 ;
        RECT 32.480 200.890 32.710 200.900 ;
        RECT 35.970 200.890 36.330 201.220 ;
        RECT 36.845 201.100 40.845 201.240 ;
        RECT 36.845 201.055 37.135 201.100 ;
        RECT 38.035 201.055 38.325 201.100 ;
        RECT 40.555 201.055 40.845 201.100 ;
        RECT 32.480 200.870 36.330 200.890 ;
        RECT 12.500 200.530 20.280 200.640 ;
        RECT 23.620 200.590 24.010 200.640 ;
        RECT 24.860 200.640 36.330 200.870 ;
        RECT 24.860 200.540 32.710 200.640 ;
        RECT 35.970 200.600 36.330 200.640 ;
        RECT 37.200 200.890 37.570 200.920 ;
        RECT 44.780 200.890 45.050 200.950 ;
        RECT 37.200 200.620 45.050 200.890 ;
        RECT 44.780 200.560 45.050 200.620 ;
        RECT 12.500 200.520 12.770 200.530 ;
        RECT 20.050 200.480 20.280 200.530 ;
        RECT 24.870 200.520 25.270 200.540 ;
        RECT 8.000 199.800 9.040 200.300 ;
        RECT 17.990 200.040 18.850 200.320 ;
        RECT 20.970 200.200 21.430 200.500 ;
        RECT 32.480 200.490 32.710 200.540 ;
        RECT 30.410 200.080 31.280 200.350 ;
        RECT 33.700 200.090 34.040 200.340 ;
        RECT 42.720 200.060 43.660 200.360 ;
        RECT 45.790 199.970 46.110 200.420 ;
        RECT 20.800 199.900 23.680 199.910 ;
        RECT 8.040 199.780 9.040 199.800 ;
        RECT 11.140 199.850 33.220 199.900 ;
        RECT 35.880 199.850 45.540 199.880 ;
        RECT 11.140 199.420 45.540 199.850 ;
        RECT 55.530 199.560 58.130 202.060 ;
        RECT 21.860 199.030 22.990 199.420 ;
        RECT 33.170 199.400 45.540 199.420 ;
        RECT 33.170 199.380 35.970 199.400 ;
        RECT 21.860 198.330 50.440 199.030 ;
        RECT 21.930 198.030 50.440 198.330 ;
        RECT 82.460 198.200 83.460 206.660 ;
        RECT 84.560 204.710 85.280 206.210 ;
        RECT 114.990 206.160 117.360 209.140 ;
        RECT 129.800 206.920 131.000 208.220 ;
        RECT 131.760 207.040 132.760 207.130 ;
        RECT 131.760 206.920 132.890 207.040 ;
        RECT 129.800 206.280 132.890 206.920 ;
        RECT 129.800 206.200 132.760 206.280 ;
        RECT 129.800 206.190 131.000 206.200 ;
        RECT 114.990 206.150 118.340 206.160 ;
        RECT 86.590 205.670 118.340 206.150 ;
        RECT 131.760 206.130 132.760 206.200 ;
        RECT 93.980 205.130 94.270 205.175 ;
        RECT 95.550 205.130 95.840 205.175 ;
        RECT 97.650 205.130 97.940 205.175 ;
        RECT 93.980 204.990 97.940 205.130 ;
        RECT 93.980 204.945 94.270 204.990 ;
        RECT 95.550 204.945 95.840 204.990 ;
        RECT 97.650 204.945 97.940 204.990 ;
        RECT 103.580 205.130 103.870 205.175 ;
        RECT 105.150 205.130 105.440 205.175 ;
        RECT 107.250 205.130 107.540 205.175 ;
        RECT 103.580 204.990 107.540 205.130 ;
        RECT 103.580 204.945 103.870 204.990 ;
        RECT 105.150 204.945 105.440 204.990 ;
        RECT 107.250 204.945 107.540 204.990 ;
        RECT 112.490 205.130 112.780 205.175 ;
        RECT 114.060 205.130 114.350 205.175 ;
        RECT 116.160 205.130 116.450 205.175 ;
        RECT 117.340 205.160 118.340 205.670 ;
        RECT 112.490 204.990 116.450 205.130 ;
        RECT 112.490 204.945 112.780 204.990 ;
        RECT 114.060 204.945 114.350 204.990 ;
        RECT 116.160 204.945 116.450 204.990 ;
        RECT 85.430 204.900 86.370 204.930 ;
        RECT 85.430 204.710 86.590 204.900 ;
        RECT 84.560 204.680 86.590 204.710 ;
        RECT 93.545 204.790 93.835 204.835 ;
        RECT 96.065 204.790 96.355 204.835 ;
        RECT 97.255 204.790 97.545 204.835 ;
        RECT 84.560 204.110 86.600 204.680 ;
        RECT 93.545 204.650 97.545 204.790 ;
        RECT 93.545 204.605 93.835 204.650 ;
        RECT 96.065 204.605 96.355 204.650 ;
        RECT 97.255 204.605 97.545 204.650 ;
        RECT 103.145 204.790 103.435 204.835 ;
        RECT 105.665 204.790 105.955 204.835 ;
        RECT 106.855 204.790 107.145 204.835 ;
        RECT 103.145 204.650 107.145 204.790 ;
        RECT 103.145 204.605 103.435 204.650 ;
        RECT 105.665 204.605 105.955 204.650 ;
        RECT 106.855 204.605 107.145 204.650 ;
        RECT 112.055 204.790 112.345 204.835 ;
        RECT 114.575 204.790 114.865 204.835 ;
        RECT 115.765 204.790 116.055 204.835 ;
        RECT 112.055 204.650 116.055 204.790 ;
        RECT 112.055 204.605 112.345 204.650 ;
        RECT 114.575 204.605 114.865 204.650 ;
        RECT 115.765 204.605 116.055 204.650 ;
        RECT 84.560 203.930 86.590 204.110 ;
        RECT 84.560 203.730 85.430 203.930 ;
        RECT 85.590 203.900 86.590 203.930 ;
        RECT 84.590 203.710 85.430 203.730 ;
        RECT 89.140 203.880 89.430 204.490 ;
        RECT 89.830 204.450 90.120 204.490 ;
        RECT 96.860 204.450 97.150 204.510 ;
        RECT 89.830 204.120 97.150 204.450 ;
        RECT 89.830 204.030 90.120 204.120 ;
        RECT 96.860 204.050 97.150 204.120 ;
        RECT 99.430 204.350 99.720 204.390 ;
        RECT 106.470 204.350 106.760 204.410 ;
        RECT 99.430 204.020 106.760 204.350 ;
        RECT 99.430 203.930 99.720 204.020 ;
        RECT 106.470 203.950 106.760 204.020 ;
        RECT 108.370 204.270 108.620 204.320 ;
        RECT 115.410 204.270 115.660 204.330 ;
        RECT 108.370 203.990 115.660 204.270 ;
        RECT 108.370 203.930 108.620 203.990 ;
        RECT 115.410 203.940 115.660 203.990 ;
        RECT 89.140 203.870 91.590 203.880 ;
        RECT 89.140 203.600 91.630 203.870 ;
        RECT 117.000 203.630 118.430 204.700 ;
        RECT 89.140 203.590 91.590 203.600 ;
        RECT 89.180 203.580 91.590 203.590 ;
        RECT 85.590 202.950 117.480 203.430 ;
        RECT 85.590 202.080 86.590 202.950 ;
        RECT 85.360 199.540 87.220 202.080 ;
        RECT 49.050 196.600 50.350 198.030 ;
        RECT 82.460 197.200 109.410 198.200 ;
        RECT 108.340 196.700 109.340 197.200 ;
        RECT 97.030 196.240 109.340 196.700 ;
        RECT 97.030 196.220 108.070 196.240 ;
        RECT 101.815 195.680 102.105 195.725 ;
        RECT 104.935 195.680 105.225 195.725 ;
        RECT 106.825 195.680 107.115 195.725 ;
        RECT 101.815 195.540 107.115 195.680 ;
        RECT 94.280 195.250 95.380 195.510 ;
        RECT 101.815 195.495 102.105 195.540 ;
        RECT 104.935 195.495 105.225 195.540 ;
        RECT 106.825 195.495 107.115 195.540 ;
        RECT 94.280 194.630 98.900 195.250 ;
        RECT 100.735 194.705 101.025 195.020 ;
        RECT 101.815 195.000 102.105 195.045 ;
        RECT 105.395 195.000 105.685 195.045 ;
        RECT 107.230 195.000 107.520 195.045 ;
        RECT 101.815 194.860 107.520 195.000 ;
        RECT 101.815 194.815 102.105 194.860 ;
        RECT 105.395 194.815 105.685 194.860 ;
        RECT 107.230 194.815 107.520 194.860 ;
        RECT 100.435 194.660 101.025 194.705 ;
        RECT 103.675 194.660 104.325 194.705 ;
        RECT 100.435 194.650 104.325 194.660 ;
        RECT 94.280 194.610 98.890 194.630 ;
        RECT 94.280 194.510 95.380 194.610 ;
        RECT 100.435 194.520 104.340 194.650 ;
        RECT 94.330 194.460 95.330 194.510 ;
        RECT 100.435 194.475 100.725 194.520 ;
        RECT 103.640 194.350 104.340 194.520 ;
        RECT 95.480 193.960 96.490 193.970 ;
        RECT 97.030 193.960 108.070 193.980 ;
        RECT 95.480 193.500 108.070 193.960 ;
        RECT 95.480 189.640 96.490 193.500 ;
        RECT 97.690 192.900 98.430 193.230 ;
        RECT 104.290 193.140 106.750 193.150 ;
        RECT 97.740 190.760 98.380 192.900 ;
        RECT 103.560 192.690 106.750 193.140 ;
        RECT 104.290 192.680 106.750 192.690 ;
        RECT 98.770 192.340 101.530 192.350 ;
        RECT 98.770 192.330 103.710 192.340 ;
        RECT 105.200 192.330 105.740 192.340 ;
        RECT 98.770 191.890 105.740 192.330 ;
        RECT 98.770 191.870 101.530 191.890 ;
        RECT 103.390 191.880 105.740 191.890 ;
        RECT 103.390 191.850 105.690 191.880 ;
        RECT 106.100 191.090 106.750 192.680 ;
        RECT 97.740 190.450 99.380 190.760 ;
        RECT 99.750 190.140 100.120 190.720 ;
        RECT 99.690 189.870 100.170 190.140 ;
        RECT 105.290 190.090 106.750 191.090 ;
        RECT 105.290 190.070 105.570 190.090 ;
        RECT 95.480 189.610 103.770 189.640 ;
        RECT 95.480 189.150 105.690 189.610 ;
        RECT 93.370 186.620 94.620 186.630 ;
        RECT 93.370 186.490 94.630 186.620 ;
        RECT 93.370 186.460 94.840 186.490 ;
        RECT 93.370 185.830 95.130 186.460 ;
        RECT 93.370 185.800 94.840 185.830 ;
        RECT 93.370 185.630 94.630 185.800 ;
        RECT 93.630 185.620 94.630 185.630 ;
        RECT 95.480 185.220 96.490 189.150 ;
        RECT 103.390 189.130 105.690 189.150 ;
        RECT 106.100 188.780 106.750 190.090 ;
        RECT 104.240 188.770 106.750 188.780 ;
        RECT 103.520 188.340 106.750 188.770 ;
        RECT 103.520 188.320 104.310 188.340 ;
        RECT 96.910 187.940 107.950 187.950 ;
        RECT 108.290 187.940 109.340 196.240 ;
        RECT 131.730 196.890 132.730 197.020 ;
        RECT 131.730 196.130 132.850 196.890 ;
        RECT 131.730 196.020 132.730 196.130 ;
        RECT 109.990 195.380 111.680 195.540 ;
        RECT 109.770 194.720 111.680 195.380 ;
        RECT 109.990 194.540 111.680 194.720 ;
        RECT 110.710 194.420 111.680 194.540 ;
        RECT 133.130 189.920 133.610 219.400 ;
        RECT 134.720 218.640 135.090 218.890 ;
        RECT 134.720 218.360 135.080 218.640 ;
        RECT 133.830 216.980 134.140 217.070 ;
        RECT 133.830 216.610 135.690 216.980 ;
        RECT 133.830 216.600 135.450 216.610 ;
        RECT 133.830 216.440 134.140 216.600 ;
        RECT 134.780 215.840 135.100 216.330 ;
        RECT 134.445 214.415 134.675 214.705 ;
        RECT 134.105 213.980 134.335 214.270 ;
        RECT 134.150 212.700 134.290 213.980 ;
        RECT 134.105 212.410 134.335 212.700 ;
        RECT 134.150 210.600 134.290 212.410 ;
        RECT 134.490 212.185 134.630 214.415 ;
        RECT 134.445 211.895 134.675 212.185 ;
        RECT 134.490 210.995 134.630 211.895 ;
        RECT 134.830 211.440 135.080 215.840 ;
        RECT 134.800 211.070 135.090 211.440 ;
        RECT 134.445 210.705 134.675 210.995 ;
        RECT 134.105 210.310 134.335 210.600 ;
        RECT 134.680 208.520 135.050 208.770 ;
        RECT 134.680 208.200 135.040 208.520 ;
        RECT 133.800 206.820 134.110 206.960 ;
        RECT 135.380 206.820 135.690 206.860 ;
        RECT 133.800 206.490 135.690 206.820 ;
        RECT 133.800 206.330 134.110 206.490 ;
        RECT 134.720 205.600 135.040 206.010 ;
        RECT 134.720 205.520 135.080 205.600 ;
        RECT 134.445 204.295 134.675 204.585 ;
        RECT 134.105 203.860 134.335 204.150 ;
        RECT 134.150 202.580 134.290 203.860 ;
        RECT 134.105 202.290 134.335 202.580 ;
        RECT 134.150 200.480 134.290 202.290 ;
        RECT 134.490 202.065 134.630 204.295 ;
        RECT 134.445 201.775 134.675 202.065 ;
        RECT 134.490 200.875 134.630 201.775 ;
        RECT 134.850 201.320 135.080 205.520 ;
        RECT 134.800 200.950 135.090 201.320 ;
        RECT 134.445 200.585 134.675 200.875 ;
        RECT 134.105 200.190 134.335 200.480 ;
        RECT 134.680 198.440 135.050 198.690 ;
        RECT 134.690 198.090 135.050 198.440 ;
        RECT 133.870 196.750 134.180 196.850 ;
        RECT 133.870 196.380 135.690 196.750 ;
        RECT 133.870 196.350 135.430 196.380 ;
        RECT 133.870 196.220 134.180 196.350 ;
        RECT 134.820 195.370 135.140 195.860 ;
        RECT 134.445 194.185 134.675 194.475 ;
        RECT 134.105 193.750 134.335 194.040 ;
        RECT 134.150 192.470 134.290 193.750 ;
        RECT 134.105 192.180 134.335 192.470 ;
        RECT 134.150 190.370 134.290 192.180 ;
        RECT 134.490 191.955 134.630 194.185 ;
        RECT 134.445 191.665 134.675 191.955 ;
        RECT 134.490 190.765 134.630 191.665 ;
        RECT 134.820 191.090 135.130 195.370 ;
        RECT 135.850 193.480 136.330 219.400 ;
        RECT 139.980 219.220 140.680 222.010 ;
        RECT 134.830 190.840 135.120 191.090 ;
        RECT 134.445 190.475 134.675 190.765 ;
        RECT 134.105 190.080 134.335 190.370 ;
        RECT 133.120 189.510 133.610 189.920 ;
        RECT 135.850 189.680 138.070 193.480 ;
        RECT 135.850 189.510 136.330 189.680 ;
        RECT 96.910 187.480 109.340 187.940 ;
        RECT 125.180 188.850 129.620 188.920 ;
        RECT 133.120 188.870 133.590 189.510 ;
        RECT 134.550 188.890 135.110 188.950 ;
        RECT 131.600 188.850 133.590 188.870 ;
        RECT 125.180 187.870 133.590 188.850 ;
        RECT 134.350 188.490 135.350 188.890 ;
        RECT 140.140 188.490 140.480 219.220 ;
        RECT 134.350 188.150 140.480 188.490 ;
        RECT 134.350 187.890 135.350 188.150 ;
        RECT 140.140 188.050 140.480 188.150 ;
        RECT 125.180 187.850 132.740 187.870 ;
        RECT 125.180 187.830 129.620 187.850 ;
        RECT 96.910 187.470 107.950 187.480 ;
        RECT 101.695 186.930 101.985 186.975 ;
        RECT 104.815 186.930 105.105 186.975 ;
        RECT 106.705 186.930 106.995 186.975 ;
        RECT 101.695 186.790 106.995 186.930 ;
        RECT 110.640 186.800 111.660 186.810 ;
        RECT 101.695 186.745 101.985 186.790 ;
        RECT 104.815 186.745 105.105 186.790 ;
        RECT 106.705 186.745 106.995 186.790 ;
        RECT 109.880 186.640 111.660 186.800 ;
        RECT 98.470 186.470 98.780 186.480 ;
        RECT 97.040 185.840 98.780 186.470 ;
        RECT 100.615 185.955 100.905 186.270 ;
        RECT 101.695 186.250 101.985 186.295 ;
        RECT 105.275 186.250 105.565 186.295 ;
        RECT 107.110 186.250 107.400 186.295 ;
        RECT 101.695 186.110 107.400 186.250 ;
        RECT 101.695 186.065 101.985 186.110 ;
        RECT 105.275 186.065 105.565 186.110 ;
        RECT 107.110 186.065 107.400 186.110 ;
        RECT 103.610 185.955 104.290 185.960 ;
        RECT 98.470 185.830 98.780 185.840 ;
        RECT 100.315 185.910 100.905 185.955 ;
        RECT 103.555 185.910 104.290 185.955 ;
        RECT 109.590 185.950 111.660 186.640 ;
        RECT 100.315 185.770 104.290 185.910 ;
        RECT 109.880 185.800 111.660 185.950 ;
        RECT 100.315 185.725 100.605 185.770 ;
        RECT 103.555 185.725 104.290 185.770 ;
        RECT 103.610 185.670 104.290 185.725 ;
        RECT 96.910 185.220 107.950 185.230 ;
        RECT 48.840 184.770 50.740 185.140 ;
        RECT 95.480 184.770 107.950 185.220 ;
        RECT 48.840 184.760 107.950 184.770 ;
        RECT 48.840 183.760 96.515 184.760 ;
        RECT 96.910 184.750 107.950 184.760 ;
        RECT 48.840 183.380 50.740 183.760 ;
        RECT 95.480 183.560 96.490 183.760 ;
        RECT 48.800 180.680 52.490 181.600 ;
        RECT 48.800 180.640 132.650 180.680 ;
        RECT 48.800 180.600 138.010 180.640 ;
        RECT 48.800 178.160 138.040 180.600 ;
        RECT 48.800 177.680 132.650 178.160 ;
        RECT 48.800 177.000 52.490 177.680 ;
        RECT 143.720 175.120 144.220 178.440 ;
        RECT 143.790 168.855 144.180 175.120 ;
        RECT 147.400 175.070 148.020 178.580 ;
        RECT 40.540 155.300 47.680 155.320 ;
        RECT 76.960 155.300 78.360 155.330 ;
        RECT 40.540 153.920 78.360 155.300 ;
        RECT 47.590 153.900 78.360 153.920 ;
        RECT 0.960 152.520 11.860 153.490 ;
        RECT 76.960 153.190 78.360 153.900 ;
        RECT 0.960 151.270 72.590 152.520 ;
        RECT 76.890 152.130 78.360 153.190 ;
        RECT 76.890 151.940 78.260 152.130 ;
        RECT 0.960 150.280 76.490 151.270 ;
        RECT 0.960 148.920 11.860 150.280 ;
        RECT 56.360 150.000 76.490 150.280 ;
        RECT 56.360 149.660 75.790 150.000 ;
        RECT 56.360 149.650 75.750 149.660 ;
        RECT 51.730 147.140 55.840 149.330 ;
        RECT 56.360 146.550 57.570 149.650 ;
        RECT 77.090 149.580 78.090 151.940 ;
        RECT 78.500 150.490 88.270 151.380 ;
        RECT 101.810 150.590 103.170 151.900 ;
        RECT 78.500 149.890 88.350 150.490 ;
        RECT 78.500 149.880 88.400 149.890 ;
        RECT 85.060 149.860 88.400 149.880 ;
        RECT 77.090 149.280 79.620 149.580 ;
        RECT 80.870 149.310 82.780 149.590 ;
        RECT 80.890 149.300 81.360 149.310 ;
        RECT 82.470 149.300 82.760 149.310 ;
        RECT 77.090 149.180 78.090 149.280 ;
        RECT 59.045 149.110 59.335 149.155 ;
        RECT 60.935 149.110 61.225 149.155 ;
        RECT 64.055 149.110 64.345 149.155 ;
        RECT 59.045 148.970 64.345 149.110 ;
        RECT 81.150 149.095 81.360 149.300 ;
        RECT 83.950 149.240 84.430 149.630 ;
        RECT 85.550 149.200 88.400 149.860 ;
        RECT 89.280 149.850 97.960 149.880 ;
        RECT 89.280 149.540 98.000 149.850 ;
        RECT 102.190 149.780 102.820 150.590 ;
        RECT 59.045 148.925 59.335 148.970 ;
        RECT 60.935 148.925 61.225 148.970 ;
        RECT 64.055 148.925 64.345 148.970 ;
        RECT 67.230 148.910 67.610 148.920 ;
        RECT 70.970 148.910 71.970 149.060 ;
        RECT 67.230 148.830 71.970 148.910 ;
        RECT 58.640 148.430 58.930 148.475 ;
        RECT 60.475 148.430 60.765 148.475 ;
        RECT 64.055 148.430 64.345 148.475 ;
        RECT 58.640 148.290 64.345 148.430 ;
        RECT 58.640 148.245 58.930 148.290 ;
        RECT 60.475 148.245 60.765 148.290 ;
        RECT 64.055 148.245 64.345 148.290 ;
        RECT 65.135 148.135 65.425 148.450 ;
        RECT 67.230 148.270 72.000 148.830 ;
        RECT 77.070 148.590 77.640 148.640 ;
        RECT 77.070 148.580 78.160 148.590 ;
        RECT 67.230 148.230 67.610 148.270 ;
        RECT 61.835 148.090 62.485 148.135 ;
        RECT 62.805 148.090 63.365 148.110 ;
        RECT 65.135 148.090 65.725 148.135 ;
        RECT 70.930 148.090 72.000 148.270 ;
        RECT 75.650 148.200 78.160 148.580 ;
        RECT 61.835 147.950 65.725 148.090 ;
        RECT 70.970 148.060 71.970 148.090 ;
        RECT 61.835 147.905 62.485 147.950 ;
        RECT 62.805 147.780 63.365 147.950 ;
        RECT 65.435 147.905 65.725 147.950 ;
        RECT 68.990 147.420 70.530 148.040 ;
        RECT 68.920 147.410 70.570 147.420 ;
        RECT 58.090 146.930 70.570 147.410 ;
        RECT 56.310 146.380 57.570 146.550 ;
        RECT 62.350 146.430 65.150 146.450 ;
        RECT 60.240 146.380 61.330 146.390 ;
        RECT 62.350 146.380 67.730 146.430 ;
        RECT 56.310 145.950 67.730 146.380 ;
        RECT 69.200 146.130 70.570 146.930 ;
        RECT 56.310 145.910 65.150 145.950 ;
        RECT 56.310 145.900 62.560 145.910 ;
        RECT 56.310 145.880 60.290 145.900 ;
        RECT 56.310 145.810 57.570 145.880 ;
        RECT 56.360 142.720 57.570 145.810 ;
        RECT 59.170 144.270 60.020 145.000 ;
        RECT 63.880 144.760 64.840 144.830 ;
        RECT 66.350 144.810 66.810 144.890 ;
        RECT 63.870 144.480 64.840 144.760 ;
        RECT 63.880 144.450 64.840 144.480 ;
        RECT 66.310 144.520 66.810 144.810 ;
        RECT 66.310 144.470 66.750 144.520 ;
        RECT 69.210 144.490 70.540 146.130 ;
        RECT 71.080 145.420 71.880 148.060 ;
        RECT 75.650 147.900 78.110 148.200 ;
        RECT 77.070 147.590 78.110 147.900 ;
        RECT 72.720 146.930 75.520 147.410 ;
        RECT 78.570 147.380 78.810 147.390 ;
        RECT 79.120 147.380 79.350 149.095 ;
        RECT 78.570 147.110 79.350 147.380 ;
        RECT 68.750 144.460 70.540 144.490 ;
        RECT 71.030 144.470 72.200 145.420 ;
        RECT 78.570 145.250 78.810 147.110 ;
        RECT 79.120 147.095 79.350 147.110 ;
        RECT 79.560 147.095 79.790 149.095 ;
        RECT 80.700 147.095 80.930 149.095 ;
        RECT 81.140 147.440 81.370 149.095 ;
        RECT 81.080 147.100 81.440 147.440 ;
        RECT 81.140 147.095 81.370 147.100 ;
        RECT 82.280 147.095 82.510 149.095 ;
        RECT 82.720 148.200 82.950 149.095 ;
        RECT 83.860 148.200 84.090 149.095 ;
        RECT 82.720 147.960 84.090 148.200 ;
        RECT 82.720 147.095 82.950 147.960 ;
        RECT 83.860 147.095 84.090 147.960 ;
        RECT 84.300 147.310 84.530 149.095 ;
        RECT 85.590 148.940 88.400 149.200 ;
        RECT 88.780 149.400 89.160 149.420 ;
        RECT 88.780 149.365 89.280 149.400 ;
        RECT 92.960 149.365 93.390 149.370 ;
        RECT 85.590 148.780 88.350 148.940 ;
        RECT 88.780 148.770 89.350 149.365 ;
        RECT 88.730 148.565 89.350 148.770 ;
        RECT 89.560 148.565 89.790 149.365 ;
        RECT 90.940 149.355 91.230 149.360 ;
        RECT 90.940 148.770 91.460 149.355 ;
        RECT 88.730 148.180 89.150 148.565 ;
        RECT 90.890 148.555 91.460 148.770 ;
        RECT 91.670 148.555 91.900 149.355 ;
        RECT 92.960 148.770 93.570 149.365 ;
        RECT 92.910 148.565 93.570 148.770 ;
        RECT 93.780 148.565 94.010 149.365 ;
        RECT 96.770 148.565 97.000 149.365 ;
        RECT 97.210 149.070 97.440 149.365 ;
        RECT 97.710 149.070 98.000 149.540 ;
        RECT 99.180 149.520 102.820 149.780 ;
        RECT 99.190 149.490 101.150 149.520 ;
        RECT 98.910 149.070 99.140 149.330 ;
        RECT 97.210 148.780 99.140 149.070 ;
        RECT 97.210 148.565 97.440 148.780 ;
        RECT 89.310 148.330 89.600 148.360 ;
        RECT 88.720 147.850 89.150 148.180 ;
        RECT 89.290 148.080 89.620 148.330 ;
        RECT 85.100 147.310 86.750 147.370 ;
        RECT 84.300 147.100 86.750 147.310 ;
        RECT 84.300 147.095 84.530 147.100 ;
        RECT 79.290 146.630 79.610 146.910 ;
        RECT 80.860 146.610 81.210 146.890 ;
        RECT 82.470 146.860 82.760 146.890 ;
        RECT 84.050 146.870 84.340 146.890 ;
        RECT 82.450 146.610 82.780 146.860 ;
        RECT 84.020 146.610 84.370 146.870 ;
        RECT 85.100 146.590 86.750 147.100 ;
        RECT 88.710 146.940 89.610 147.850 ;
        RECT 90.890 147.840 91.230 148.555 ;
        RECT 91.420 148.320 91.710 148.350 ;
        RECT 91.400 148.070 91.730 148.320 ;
        RECT 90.740 147.080 91.630 147.840 ;
        RECT 92.910 146.750 93.350 148.565 ;
        RECT 98.910 148.530 99.140 148.780 ;
        RECT 101.200 148.530 101.430 149.330 ;
        RECT 93.530 148.330 93.820 148.360 ;
        RECT 96.960 148.330 97.250 148.360 ;
        RECT 99.190 148.350 101.150 148.370 ;
        RECT 102.190 148.350 102.820 149.520 ;
        RECT 103.580 148.900 104.600 150.500 ;
        RECT 93.510 148.080 93.840 148.330 ;
        RECT 96.940 148.080 97.270 148.330 ;
        RECT 99.170 148.090 102.820 148.350 ;
        RECT 85.090 146.300 86.750 146.590 ;
        RECT 78.570 144.980 83.180 145.250 ;
        RECT 84.550 145.010 84.890 145.270 ;
        RECT 84.575 144.980 84.865 145.010 ;
        RECT 79.740 144.820 79.910 144.980 ;
        RECT 85.100 144.910 86.750 146.300 ;
        RECT 88.380 146.560 88.630 146.580 ;
        RECT 88.380 146.270 88.660 146.560 ;
        RECT 88.865 146.520 98.865 146.750 ;
        RECT 99.090 146.560 99.360 146.590 ;
        RECT 88.380 146.250 88.630 146.270 ;
        RECT 88.865 146.080 98.865 146.310 ;
        RECT 99.070 146.270 99.360 146.560 ;
        RECT 93.980 145.230 94.950 146.080 ;
        RECT 99.090 145.570 99.360 146.270 ;
        RECT 88.320 145.220 94.950 145.230 ;
        RECT 85.100 144.820 85.290 144.910 ;
        RECT 77.100 144.740 78.190 144.810 ;
        RECT 65.365 143.710 65.735 143.720 ;
        RECT 67.670 143.710 70.540 144.460 ;
        RECT 62.470 143.660 70.540 143.710 ;
        RECT 60.260 143.180 70.540 143.660 ;
        RECT 71.390 143.620 72.390 143.650 ;
        RECT 77.090 143.620 78.190 144.740 ;
        RECT 79.120 143.820 79.350 144.820 ;
        RECT 79.710 143.820 79.940 144.820 ;
        RECT 80.850 143.820 81.080 144.820 ;
        RECT 81.440 144.810 81.670 144.820 ;
        RECT 81.390 144.470 81.750 144.810 ;
        RECT 81.440 143.820 81.670 144.470 ;
        RECT 82.580 143.820 82.810 144.820 ;
        RECT 83.170 144.310 83.400 144.820 ;
        RECT 84.310 144.310 84.540 144.820 ;
        RECT 83.170 144.090 84.540 144.310 ;
        RECT 83.170 143.820 83.400 144.090 ;
        RECT 84.310 143.820 84.540 144.090 ;
        RECT 84.900 144.570 85.290 144.820 ;
        RECT 88.300 144.860 94.950 145.220 ;
        RECT 98.180 145.020 99.460 145.570 ;
        RECT 102.190 145.480 102.820 148.090 ;
        RECT 103.610 146.200 104.570 148.900 ;
        RECT 100.970 145.250 102.930 145.480 ;
        RECT 100.550 145.130 100.760 145.150 ;
        RECT 100.530 145.090 100.760 145.130 ;
        RECT 84.900 143.820 85.130 144.570 ;
        RECT 85.800 143.755 86.800 143.770 ;
        RECT 79.385 143.650 79.675 143.660 ;
        RECT 81.115 143.650 81.405 143.660 ;
        RECT 82.845 143.650 83.135 143.660 ;
        RECT 71.270 143.510 78.190 143.620 ;
        RECT 71.240 143.430 78.190 143.510 ;
        RECT 62.470 143.170 70.540 143.180 ;
        RECT 68.750 142.720 68.900 142.740 ;
        RECT 56.360 142.250 68.900 142.720 ;
        RECT 53.660 141.675 55.660 141.710 ;
        RECT 53.645 140.665 55.660 141.675 ;
        RECT 53.660 138.260 55.660 140.665 ;
        RECT 53.870 138.240 55.660 138.260 ;
        RECT 56.360 138.750 57.570 142.250 ;
        RECT 57.860 142.240 68.900 142.250 ;
        RECT 58.815 141.700 59.105 141.745 ;
        RECT 60.705 141.700 60.995 141.745 ;
        RECT 63.825 141.700 64.115 141.745 ;
        RECT 58.815 141.560 64.115 141.700 ;
        RECT 58.815 141.515 59.105 141.560 ;
        RECT 60.705 141.515 60.995 141.560 ;
        RECT 63.825 141.515 64.115 141.560 ;
        RECT 67.000 141.420 67.350 141.480 ;
        RECT 58.410 141.020 58.700 141.065 ;
        RECT 60.245 141.020 60.535 141.065 ;
        RECT 63.825 141.020 64.115 141.065 ;
        RECT 58.410 140.880 64.115 141.020 ;
        RECT 58.410 140.835 58.700 140.880 ;
        RECT 60.245 140.835 60.535 140.880 ;
        RECT 63.825 140.835 64.115 140.880 ;
        RECT 64.905 140.725 65.195 141.040 ;
        RECT 67.000 140.790 69.030 141.420 ;
        RECT 69.210 140.900 70.540 143.170 ;
        RECT 70.840 142.680 78.190 143.430 ;
        RECT 79.350 143.380 83.170 143.650 ;
        RECT 84.480 143.340 84.950 143.660 ;
        RECT 71.270 142.620 78.190 142.680 ;
        RECT 77.100 142.610 78.190 142.620 ;
        RECT 85.455 142.770 86.800 143.755 ;
        RECT 84.000 142.015 85.130 142.020 ;
        RECT 85.455 142.015 86.785 142.770 ;
        RECT 88.300 142.370 88.630 144.860 ;
        RECT 93.980 144.640 94.950 144.860 ;
        RECT 93.480 144.450 93.730 144.470 ;
        RECT 93.480 144.160 93.760 144.450 ;
        RECT 93.920 144.410 98.920 144.640 ;
        RECT 99.090 144.450 99.360 145.020 ;
        RECT 93.480 144.140 93.730 144.160 ;
        RECT 93.920 143.990 98.920 144.200 ;
        RECT 99.080 144.160 99.360 144.450 ;
        RECT 99.090 144.140 99.360 144.160 ;
        RECT 100.530 144.290 100.920 145.090 ;
        RECT 100.530 143.990 100.760 144.290 ;
        RECT 102.190 144.130 102.820 145.250 ;
        RECT 102.980 144.290 103.210 145.090 ;
        RECT 93.920 143.980 99.980 143.990 ;
        RECT 100.160 143.980 100.760 143.990 ;
        RECT 93.920 143.970 100.760 143.980 ;
        RECT 97.970 143.770 100.760 143.970 ;
        RECT 100.970 143.900 102.930 144.130 ;
        RECT 97.970 143.760 100.750 143.770 ;
        RECT 90.180 142.510 91.870 142.670 ;
        RECT 88.260 142.350 88.630 142.370 ;
        RECT 69.210 140.850 70.550 140.900 ;
        RECT 84.000 140.885 86.795 142.015 ;
        RECT 88.260 141.110 88.700 142.350 ;
        RECT 88.855 142.280 98.855 142.510 ;
        RECT 99.080 142.320 99.350 142.350 ;
        RECT 88.855 141.840 98.855 142.070 ;
        RECT 99.060 142.030 99.350 142.320 ;
        RECT 88.260 141.090 88.670 141.110 ;
        RECT 93.970 141.010 95.370 141.840 ;
        RECT 99.080 141.560 99.350 142.030 ;
        RECT 98.350 141.110 99.390 141.560 ;
        RECT 102.190 141.240 102.820 143.900 ;
        RECT 84.000 140.850 85.130 140.885 ;
        RECT 61.605 140.680 62.255 140.725 ;
        RECT 63.210 140.680 63.760 140.690 ;
        RECT 64.905 140.680 65.495 140.725 ;
        RECT 67.000 140.720 67.350 140.790 ;
        RECT 69.210 140.700 85.130 140.850 ;
        RECT 61.605 140.540 65.495 140.680 ;
        RECT 61.605 140.495 62.255 140.540 ;
        RECT 63.210 140.420 63.760 140.540 ;
        RECT 65.205 140.495 65.495 140.540 ;
        RECT 69.170 140.010 85.130 140.700 ;
        RECT 91.240 140.570 95.370 141.010 ;
        RECT 68.830 140.000 85.130 140.010 ;
        RECT 57.860 139.520 85.130 140.000 ;
        RECT 91.200 140.540 95.370 140.570 ;
        RECT 91.200 139.830 92.370 140.540 ;
        RECT 93.970 140.390 95.370 140.540 ;
        RECT 93.460 140.200 93.710 140.220 ;
        RECT 93.460 139.910 93.740 140.200 ;
        RECT 93.900 140.160 98.900 140.390 ;
        RECT 99.080 140.200 99.350 141.110 ;
        RECT 100.950 141.010 102.910 141.240 ;
        RECT 100.670 140.840 100.900 140.850 ;
        RECT 100.370 140.300 100.900 140.840 ;
        RECT 93.460 139.890 93.710 139.910 ;
        RECT 88.640 139.800 92.370 139.830 ;
        RECT 71.430 138.750 83.290 138.760 ;
        RECT 56.360 138.300 83.290 138.750 ;
        RECT 54.155 129.810 55.165 138.240 ;
        RECT 56.360 135.220 57.570 138.300 ;
        RECT 71.430 138.280 83.290 138.300 ;
        RECT 76.560 137.740 76.850 137.785 ;
        RECT 78.130 137.740 78.420 137.785 ;
        RECT 80.230 137.740 80.520 137.785 ;
        RECT 76.560 137.600 80.520 137.740 ;
        RECT 76.560 137.555 76.850 137.600 ;
        RECT 78.130 137.555 78.420 137.600 ;
        RECT 80.230 137.555 80.520 137.600 ;
        RECT 71.990 137.280 72.300 137.530 ;
        RECT 72.000 137.060 72.300 137.280 ;
        RECT 76.125 137.400 76.415 137.445 ;
        RECT 78.645 137.400 78.935 137.445 ;
        RECT 79.835 137.400 80.125 137.445 ;
        RECT 76.125 137.260 80.125 137.400 ;
        RECT 76.125 137.215 76.415 137.260 ;
        RECT 78.645 137.215 78.935 137.260 ;
        RECT 79.835 137.215 80.125 137.260 ;
        RECT 79.490 137.060 79.780 137.080 ;
        RECT 69.540 135.900 70.540 136.900 ;
        RECT 72.000 136.790 79.780 137.060 ;
        RECT 72.000 136.780 79.760 136.790 ;
        RECT 79.350 136.770 79.490 136.780 ;
        RECT 73.840 136.200 74.250 136.500 ;
        RECT 71.430 135.560 81.090 136.040 ;
        RECT 71.410 135.220 81.070 135.240 ;
        RECT 81.690 135.220 81.890 138.280 ;
        RECT 82.290 137.760 83.290 138.280 ;
        RECT 82.270 137.110 83.270 137.120 ;
        RECT 56.360 135.190 81.070 135.220 ;
        RECT 81.670 135.190 81.890 135.220 ;
        RECT 56.360 134.790 81.890 135.190 ;
        RECT 82.230 134.900 83.360 137.110 ;
        RECT 56.360 134.770 81.070 134.790 ;
        RECT 56.360 131.720 57.570 134.770 ;
        RECT 71.410 134.760 81.070 134.770 ;
        RECT 76.540 134.220 76.830 134.265 ;
        RECT 78.110 134.220 78.400 134.265 ;
        RECT 80.210 134.220 80.500 134.265 ;
        RECT 76.540 134.080 80.500 134.220 ;
        RECT 71.950 133.780 72.290 134.040 ;
        RECT 76.540 134.035 76.830 134.080 ;
        RECT 78.110 134.035 78.400 134.080 ;
        RECT 80.210 134.035 80.500 134.080 ;
        RECT 76.105 133.880 76.395 133.925 ;
        RECT 78.625 133.880 78.915 133.925 ;
        RECT 79.815 133.880 80.105 133.925 ;
        RECT 71.960 133.540 72.220 133.780 ;
        RECT 76.105 133.740 80.105 133.880 ;
        RECT 76.105 133.695 76.395 133.740 ;
        RECT 78.625 133.695 78.915 133.740 ;
        RECT 79.815 133.695 80.105 133.740 ;
        RECT 80.670 133.580 81.090 133.600 ;
        RECT 79.430 133.540 79.700 133.560 ;
        RECT 71.950 133.500 79.700 133.540 ;
        RECT 71.950 133.330 79.770 133.500 ;
        RECT 69.490 132.320 70.490 133.320 ;
        RECT 72.690 133.240 79.770 133.330 ;
        RECT 80.630 133.240 81.090 133.580 ;
        RECT 72.690 133.200 79.750 133.240 ;
        RECT 73.800 132.670 74.190 132.960 ;
        RECT 71.410 132.040 81.070 132.520 ;
        RECT 71.470 131.720 81.130 131.730 ;
        RECT 56.360 131.670 81.130 131.720 ;
        RECT 81.670 131.680 81.890 134.790 ;
        RECT 84.000 134.670 85.130 139.520 ;
        RECT 88.190 139.220 92.370 139.800 ;
        RECT 93.900 139.740 98.900 139.950 ;
        RECT 99.060 139.910 99.350 140.200 ;
        RECT 100.310 140.120 100.900 140.300 ;
        RECT 99.080 139.880 99.350 139.910 ;
        RECT 100.370 140.050 100.900 140.120 ;
        RECT 99.940 139.740 100.120 139.800 ;
        RECT 100.370 139.740 100.760 140.050 ;
        RECT 102.190 139.890 102.820 141.010 ;
        RECT 102.960 140.050 103.190 140.850 ;
        RECT 93.900 139.720 100.760 139.740 ;
        RECT 98.090 139.430 100.760 139.720 ;
        RECT 100.950 139.660 102.910 139.890 ;
        RECT 98.690 139.410 100.130 139.430 ;
        RECT 100.370 139.420 100.760 139.430 ;
        RECT 88.190 138.090 88.630 139.220 ;
        RECT 91.200 139.170 92.370 139.220 ;
        RECT 97.790 138.640 99.360 139.240 ;
        RECT 88.800 138.280 92.200 138.490 ;
        RECT 88.190 137.800 88.650 138.090 ;
        RECT 88.800 138.050 98.855 138.280 ;
        RECT 99.040 138.120 99.330 138.640 ;
        RECT 88.800 138.040 92.200 138.050 ;
        RECT 88.190 137.780 88.630 137.800 ;
        RECT 88.855 137.610 98.855 137.840 ;
        RECT 93.980 137.410 94.920 137.610 ;
        RECT 99.040 137.500 99.350 138.120 ;
        RECT 91.330 137.180 94.920 137.410 ;
        RECT 88.250 135.250 89.360 136.320 ;
        RECT 89.720 135.310 90.200 136.690 ;
        RECT 91.330 136.600 91.580 137.180 ;
        RECT 93.980 137.090 94.920 137.180 ;
        RECT 93.990 136.700 94.920 137.090 ;
        RECT 91.320 136.330 91.650 136.600 ;
        RECT 92.440 135.310 92.920 136.690 ;
        RECT 93.980 136.160 94.920 136.700 ;
        RECT 93.470 135.970 93.720 135.990 ;
        RECT 93.470 135.680 93.750 135.970 ;
        RECT 93.910 135.930 98.910 136.160 ;
        RECT 99.090 135.970 99.350 137.500 ;
        RECT 102.190 137.000 102.820 139.660 ;
        RECT 100.960 136.770 102.920 137.000 ;
        RECT 93.470 135.660 93.720 135.680 ;
        RECT 93.910 135.520 98.910 135.720 ;
        RECT 99.070 135.680 99.350 135.970 ;
        RECT 99.090 135.660 99.350 135.680 ;
        RECT 100.420 136.610 100.820 136.630 ;
        RECT 100.420 135.810 100.910 136.610 ;
        RECT 100.420 135.520 100.820 135.810 ;
        RECT 102.190 135.650 102.820 136.770 ;
        RECT 102.970 135.810 103.200 136.610 ;
        RECT 103.590 135.860 104.590 146.200 ;
        RECT 93.910 135.490 100.820 135.520 ;
        RECT 97.500 135.170 100.820 135.490 ;
        RECT 100.960 135.420 102.920 135.650 ;
        RECT 103.560 134.930 104.590 135.860 ;
        RECT 103.560 134.860 104.580 134.930 ;
        RECT 82.170 134.485 85.130 134.670 ;
        RECT 103.570 134.485 104.580 134.860 ;
        RECT 110.970 134.550 114.410 134.580 ;
        RECT 110.970 134.485 114.420 134.550 ;
        RECT 82.170 132.020 114.420 134.485 ;
        RECT 82.170 131.780 114.410 132.020 ;
        RECT 82.170 131.730 112.950 131.780 ;
        RECT 81.670 131.670 81.880 131.680 ;
        RECT 82.170 131.670 84.530 131.730 ;
        RECT 89.210 131.700 110.910 131.730 ;
        RECT 56.360 131.270 81.880 131.670 ;
        RECT 56.360 131.260 57.570 131.270 ;
        RECT 71.470 131.250 81.130 131.270 ;
        RECT 76.600 130.710 76.890 130.755 ;
        RECT 78.170 130.710 78.460 130.755 ;
        RECT 80.270 130.710 80.560 130.755 ;
        RECT 76.600 130.570 80.560 130.710 ;
        RECT 71.990 130.260 72.340 130.530 ;
        RECT 76.600 130.525 76.890 130.570 ;
        RECT 78.170 130.525 78.460 130.570 ;
        RECT 80.270 130.525 80.560 130.570 ;
        RECT 76.165 130.370 76.455 130.415 ;
        RECT 78.685 130.370 78.975 130.415 ;
        RECT 79.875 130.370 80.165 130.415 ;
        RECT 72.050 130.000 72.280 130.260 ;
        RECT 76.165 130.230 80.165 130.370 ;
        RECT 76.165 130.185 76.455 130.230 ;
        RECT 78.685 130.185 78.975 130.230 ;
        RECT 79.875 130.185 80.165 130.230 ;
        RECT 80.690 130.070 81.130 130.080 ;
        RECT 79.450 130.010 79.780 130.020 ;
        RECT 72.890 130.000 79.790 130.010 ;
        RECT 54.155 129.800 70.270 129.810 ;
        RECT 54.155 128.800 70.440 129.800 ;
        RECT 72.040 129.760 79.790 130.000 ;
        RECT 72.890 129.750 79.790 129.760 ;
        RECT 80.660 129.740 81.130 130.070 ;
        RECT 73.890 129.420 74.240 129.450 ;
        RECT 73.870 129.160 74.290 129.420 ;
        RECT 71.470 128.530 81.130 129.010 ;
        RECT 81.360 128.560 83.600 131.090 ;
        RECT 85.170 129.770 87.620 131.270 ;
        RECT 108.720 129.780 111.090 131.320 ;
        RECT 111.450 129.100 112.950 131.730 ;
        RECT 82.270 128.540 83.280 128.560 ;
        RECT 111.595 125.485 112.925 129.100 ;
        RECT 143.830 33.360 144.130 168.855 ;
        RECT 113.050 31.700 118.240 33.150 ;
        RECT 115.030 30.520 116.420 31.700 ;
        RECT 114.920 29.630 116.420 30.520 ;
        RECT 143.690 30.370 144.280 33.360 ;
        RECT 147.515 32.720 147.815 175.070 ;
        RECT 147.300 30.310 148.060 32.720 ;
        RECT 114.920 29.520 115.920 29.630 ;
        RECT 115.060 29.380 115.840 29.520 ;
        RECT 115.030 28.640 115.880 29.380 ;
        RECT 144.440 28.660 145.740 29.890 ;
        RECT 125.260 28.040 125.620 28.050 ;
        RECT 107.080 27.950 125.620 28.040 ;
        RECT 107.070 27.720 125.620 27.950 ;
        RECT 143.170 27.790 145.270 28.440 ;
        RECT 151.840 28.030 153.000 29.590 ;
        RECT 107.080 27.670 125.620 27.720 ;
        RECT 106.190 27.510 106.540 27.570 ;
        RECT 106.170 26.860 106.560 27.510 ;
        RECT 106.790 27.450 107.020 27.515 ;
        RECT 106.190 26.800 106.540 26.860 ;
        RECT 106.740 26.820 107.100 27.450 ;
        RECT 106.790 24.265 107.020 26.820 ;
        RECT 107.880 24.870 108.110 27.515 ;
        RECT 108.970 27.470 109.200 27.515 ;
        RECT 111.910 27.480 112.140 27.515 ;
        RECT 108.960 26.840 109.320 27.470 ;
        RECT 111.290 27.400 111.640 27.460 ;
        RECT 107.800 24.320 108.190 24.870 ;
        RECT 107.880 24.265 108.110 24.320 ;
        RECT 108.970 24.265 109.200 26.840 ;
        RECT 111.270 26.700 111.660 27.400 ;
        RECT 111.800 26.780 112.190 27.480 ;
        RECT 111.290 26.640 111.640 26.700 ;
        RECT 111.910 24.265 112.140 26.780 ;
        RECT 113.000 24.940 113.230 27.515 ;
        RECT 114.090 27.440 114.320 27.515 ;
        RECT 114.060 26.740 114.450 27.440 ;
        RECT 112.920 24.310 113.300 24.940 ;
        RECT 113.000 24.265 113.230 24.310 ;
        RECT 114.090 24.265 114.320 26.740 ;
        RECT 116.350 26.710 116.750 27.500 ;
        RECT 117.030 27.480 117.260 27.505 ;
        RECT 116.950 26.850 117.310 27.480 ;
        RECT 117.030 24.255 117.260 26.850 ;
        RECT 118.120 25.070 118.350 27.505 ;
        RECT 119.210 27.440 119.440 27.505 ;
        RECT 119.140 26.810 119.500 27.440 ;
        RECT 118.030 24.280 118.430 25.070 ;
        RECT 118.120 24.255 118.350 24.280 ;
        RECT 119.210 24.255 119.440 26.810 ;
        RECT 121.480 26.760 121.890 27.530 ;
        RECT 122.090 26.880 122.450 27.510 ;
        RECT 123.220 26.890 123.500 27.670 ;
        RECT 122.150 24.255 122.380 26.880 ;
        RECT 123.240 24.970 123.470 26.890 ;
        RECT 124.280 26.880 124.640 27.510 ;
        RECT 123.160 24.270 123.550 24.970 ;
        RECT 123.240 24.255 123.470 24.270 ;
        RECT 124.330 24.255 124.560 26.880 ;
        RECT 125.260 24.110 125.620 27.670 ;
        RECT 151.865 27.330 152.155 27.340 ;
        RECT 152.455 27.330 152.745 27.340 ;
        RECT 150.670 27.310 152.745 27.330 ;
        RECT 138.420 27.250 141.370 27.280 ;
        RECT 138.070 26.900 141.370 27.250 ;
        RECT 150.670 27.140 153.130 27.310 ;
        RECT 138.070 24.480 138.840 26.900 ;
        RECT 139.835 26.880 140.125 26.900 ;
        RECT 140.425 26.880 140.715 26.900 ;
        RECT 141.015 26.880 141.305 26.900 ;
        RECT 146.940 26.820 147.340 26.850 ;
        RECT 107.050 23.740 125.620 24.110 ;
        RECT 125.260 23.730 125.620 23.740 ;
        RECT 103.680 23.060 104.190 23.150 ;
        RECT 109.660 23.060 110.190 23.070 ;
        RECT 103.680 22.760 116.270 23.060 ;
        RECT 136.790 23.010 138.840 24.480 ;
        RECT 103.830 22.740 116.270 22.760 ;
        RECT 102.180 22.510 102.510 22.530 ;
        RECT 120.020 22.520 120.890 22.540 ;
        RECT 114.680 22.510 120.890 22.520 ;
        RECT 102.180 22.500 103.080 22.510 ;
        RECT 108.790 22.500 120.890 22.510 ;
        RECT 102.180 22.200 120.890 22.500 ;
        RECT 102.180 22.190 120.210 22.200 ;
        RECT 102.180 21.340 102.510 22.190 ;
        RECT 103.040 22.180 120.210 22.190 ;
        RECT 103.040 22.170 114.680 22.180 ;
        RECT 103.040 22.150 108.830 22.170 ;
        RECT 100.620 21.330 102.510 21.340 ;
        RECT 100.620 21.040 102.520 21.330 ;
        RECT 104.620 21.260 108.460 21.270 ;
        RECT 120.530 21.260 120.870 22.200 ;
        RECT 125.120 21.960 125.530 21.970 ;
        RECT 122.340 21.630 125.530 21.960 ;
        RECT 104.620 21.240 108.790 21.260 ;
        RECT 110.680 21.240 114.850 21.260 ;
        RECT 99.270 20.860 99.650 20.920 ;
        RECT 99.250 20.430 99.670 20.860 ;
        RECT 99.270 20.370 99.650 20.430 ;
        RECT 99.940 19.370 100.170 20.865 ;
        RECT 100.420 20.860 100.650 20.865 ;
        RECT 100.330 20.430 100.750 20.860 ;
        RECT 99.870 18.950 100.230 19.370 ;
        RECT 99.940 18.865 100.170 18.950 ;
        RECT 100.420 18.865 100.650 20.430 ;
        RECT 100.900 19.340 101.130 20.865 ;
        RECT 101.280 20.440 101.700 20.870 ;
        RECT 100.840 18.920 101.200 19.340 ;
        RECT 100.900 18.865 101.130 18.920 ;
        RECT 101.380 18.865 101.610 20.440 ;
        RECT 102.180 19.100 102.520 21.040 ;
        RECT 104.610 21.010 108.790 21.240 ;
        RECT 110.670 21.010 114.850 21.240 ;
        RECT 104.620 21.000 108.790 21.010 ;
        RECT 103.750 20.840 104.010 20.890 ;
        RECT 103.690 20.370 104.050 20.840 ;
        RECT 103.750 20.340 104.010 20.370 ;
        RECT 104.330 19.230 104.560 20.805 ;
        RECT 105.270 20.390 105.690 20.820 ;
        RECT 102.180 18.700 102.530 19.100 ;
        RECT 104.220 18.790 104.620 19.230 ;
        RECT 105.370 18.805 105.600 20.390 ;
        RECT 106.410 19.260 106.640 20.805 ;
        RECT 107.450 20.790 107.680 20.805 ;
        RECT 107.370 20.360 107.790 20.790 ;
        RECT 106.340 18.820 106.740 19.260 ;
        RECT 106.410 18.805 106.640 18.820 ;
        RECT 107.450 18.805 107.680 20.360 ;
        RECT 100.160 18.660 102.530 18.700 ;
        RECT 100.150 18.430 102.530 18.660 ;
        RECT 108.460 18.610 108.790 21.000 ;
        RECT 110.680 20.990 114.850 21.010 ;
        RECT 116.700 20.990 120.870 21.260 ;
        RECT 109.780 20.790 110.110 20.850 ;
        RECT 109.760 20.380 110.130 20.790 ;
        RECT 109.780 20.320 110.110 20.380 ;
        RECT 110.390 19.290 110.620 20.805 ;
        RECT 111.370 20.400 111.740 20.810 ;
        RECT 110.310 18.830 110.690 19.290 ;
        RECT 110.390 18.805 110.620 18.830 ;
        RECT 111.430 18.805 111.660 20.400 ;
        RECT 112.470 19.250 112.700 20.805 ;
        RECT 113.510 20.800 113.740 20.805 ;
        RECT 113.440 20.390 113.810 20.800 ;
        RECT 112.390 18.790 112.770 19.250 ;
        RECT 113.510 18.805 113.740 20.390 ;
        RECT 104.620 18.600 108.790 18.610 ;
        RECT 114.520 18.600 114.850 20.990 ;
        RECT 120.530 20.910 120.870 20.990 ;
        RECT 115.820 20.770 116.140 20.830 ;
        RECT 115.800 20.230 116.160 20.770 ;
        RECT 115.820 20.170 116.140 20.230 ;
        RECT 116.450 19.310 116.680 20.795 ;
        RECT 117.490 20.790 117.720 20.795 ;
        RECT 117.440 20.250 117.800 20.790 ;
        RECT 116.370 18.810 116.730 19.310 ;
        RECT 116.450 18.795 116.680 18.810 ;
        RECT 117.490 18.795 117.720 20.250 ;
        RECT 118.530 19.310 118.760 20.795 ;
        RECT 119.570 20.760 119.800 20.795 ;
        RECT 119.500 20.220 119.860 20.760 ;
        RECT 118.450 18.810 118.810 19.310 ;
        RECT 118.530 18.795 118.760 18.810 ;
        RECT 119.570 18.795 119.800 20.220 ;
        RECT 120.540 18.600 120.870 20.910 ;
        RECT 121.480 19.090 121.820 19.150 ;
        RECT 100.160 18.400 102.530 18.430 ;
        RECT 102.180 18.380 102.530 18.400 ;
        RECT 96.580 17.810 98.930 18.150 ;
        RECT 100.670 17.810 101.170 17.830 ;
        RECT 96.580 17.350 101.170 17.810 ;
        RECT 102.190 17.680 102.530 18.380 ;
        RECT 104.610 18.370 108.790 18.600 ;
        RECT 110.670 18.370 114.850 18.600 ;
        RECT 104.620 18.340 108.790 18.370 ;
        RECT 96.580 17.310 101.080 17.350 ;
        RECT 96.580 17.060 98.930 17.310 ;
        RECT 102.150 17.300 102.580 17.680 ;
        RECT 108.460 17.620 108.790 18.340 ;
        RECT 110.680 18.330 114.850 18.370 ;
        RECT 116.700 18.330 120.870 18.600 ;
        RECT 114.520 17.660 114.850 18.330 ;
        RECT 108.460 17.610 112.500 17.620 ;
        RECT 108.460 17.340 112.560 17.610 ;
        RECT 114.480 17.360 114.920 17.660 ;
        RECT 97.770 17.020 98.770 17.060 ;
        RECT 102.190 16.540 102.530 17.300 ;
        RECT 108.460 16.620 108.790 17.340 ;
        RECT 112.140 17.330 112.560 17.340 ;
        RECT 105.400 16.580 108.790 16.620 ;
        RECT 114.520 16.610 114.850 17.360 ;
        RECT 120.540 16.610 120.870 18.330 ;
        RECT 121.460 18.320 121.840 19.090 ;
        RECT 122.110 19.060 122.340 21.490 ;
        RECT 123.200 21.470 123.430 21.490 ;
        RECT 123.140 20.900 123.500 21.470 ;
        RECT 121.980 18.350 122.430 19.060 ;
        RECT 121.480 18.260 121.820 18.320 ;
        RECT 122.110 18.240 122.340 18.350 ;
        RECT 123.200 18.240 123.430 20.900 ;
        RECT 124.290 19.000 124.520 21.490 ;
        RECT 125.120 19.740 125.530 21.630 ;
        RECT 138.070 20.490 138.840 23.010 ;
        RECT 139.570 22.400 139.800 26.675 ;
        RECT 140.160 26.320 140.390 26.675 ;
        RECT 140.030 25.040 140.530 26.320 ;
        RECT 139.400 20.920 139.980 22.400 ;
        RECT 139.570 20.675 139.800 20.920 ;
        RECT 140.160 20.675 140.390 25.040 ;
        RECT 140.750 22.370 140.980 26.675 ;
        RECT 141.340 26.310 141.570 26.675 ;
        RECT 145.560 26.520 147.340 26.820 ;
        RECT 141.190 25.030 141.690 26.310 ;
        RECT 140.620 20.890 141.200 22.370 ;
        RECT 140.750 20.675 140.980 20.890 ;
        RECT 141.340 20.675 141.570 25.030 ;
        RECT 145.320 21.350 145.550 26.355 ;
        RECT 145.910 26.130 146.140 26.355 ;
        RECT 145.790 25.520 146.330 26.130 ;
        RECT 146.940 26.120 147.340 26.520 ;
        RECT 150.670 26.120 151.030 27.140 ;
        RECT 151.865 27.110 152.155 27.140 ;
        RECT 152.455 27.110 152.745 27.140 ;
        RECT 144.420 20.640 145.560 21.350 ;
        RECT 138.070 20.470 141.220 20.490 ;
        RECT 138.070 20.240 141.305 20.470 ;
        RECT 144.420 20.355 145.550 20.640 ;
        RECT 145.910 20.355 146.140 25.520 ;
        RECT 146.940 24.490 147.290 26.120 ;
        RECT 150.680 24.490 151.030 26.120 ;
        RECT 146.940 21.560 151.030 24.490 ;
        RECT 146.940 21.430 147.350 21.560 ;
        RECT 126.820 19.740 128.480 20.240 ;
        RECT 138.130 20.140 141.220 20.240 ;
        RECT 124.170 18.290 124.620 19.000 ;
        RECT 125.120 18.750 128.480 19.740 ;
        RECT 124.290 18.240 124.520 18.290 ;
        RECT 125.120 18.100 125.530 18.750 ;
        RECT 122.390 17.770 125.530 18.100 ;
        RECT 125.120 17.760 125.530 17.770 ;
        RECT 125.900 18.510 128.480 18.750 ;
        RECT 141.580 19.190 142.350 19.290 ;
        RECT 144.420 19.210 145.350 20.355 ;
        RECT 146.940 20.170 147.320 21.430 ;
        RECT 145.590 20.150 147.320 20.170 ;
        RECT 145.585 19.920 147.320 20.150 ;
        RECT 145.590 19.900 147.320 19.920 ;
        RECT 145.590 19.870 147.210 19.900 ;
        RECT 148.210 19.800 149.750 21.560 ;
        RECT 150.740 19.930 151.030 21.560 ;
        RECT 151.600 21.420 151.830 26.905 ;
        RECT 152.190 26.420 152.420 26.905 ;
        RECT 152.110 25.320 152.550 26.420 ;
        RECT 151.550 20.370 152.020 21.420 ;
        RECT 150.710 19.800 151.030 19.930 ;
        RECT 151.600 19.905 151.830 20.370 ;
        RECT 152.190 19.905 152.420 25.320 ;
        RECT 152.780 21.400 153.010 26.905 ;
        RECT 152.700 20.350 153.170 21.400 ;
        RECT 152.780 19.905 153.010 20.350 ;
        RECT 148.210 19.740 149.770 19.800 ;
        RECT 148.230 19.210 149.770 19.740 ;
        RECT 150.670 19.690 151.030 19.800 ;
        RECT 151.865 19.690 152.155 19.700 ;
        RECT 152.455 19.690 152.745 19.700 ;
        RECT 150.670 19.390 152.860 19.690 ;
        RECT 144.420 19.190 149.770 19.210 ;
        RECT 141.580 18.560 149.770 19.190 ;
        RECT 144.420 18.530 145.350 18.560 ;
        RECT 100.520 16.300 102.530 16.540 ;
        RECT 105.390 16.350 108.790 16.580 ;
        RECT 100.520 16.280 102.030 16.300 ;
        RECT 99.700 14.440 100.030 14.500 ;
        RECT 99.680 13.920 100.050 14.440 ;
        RECT 100.310 14.410 100.540 16.120 ;
        RECT 100.790 16.100 101.020 16.120 ;
        RECT 100.740 15.540 101.100 16.100 ;
        RECT 99.700 13.860 100.030 13.920 ;
        RECT 100.230 13.890 100.600 14.410 ;
        RECT 100.310 13.870 100.540 13.890 ;
        RECT 100.790 13.870 101.020 15.540 ;
        RECT 101.270 14.420 101.500 16.120 ;
        RECT 101.190 13.900 101.560 14.420 ;
        RECT 101.270 13.870 101.500 13.900 ;
        RECT 102.190 13.730 102.530 16.300 ;
        RECT 101.000 13.430 102.530 13.730 ;
        RECT 103.700 14.640 104.120 14.650 ;
        RECT 104.520 14.640 104.770 14.660 ;
        RECT 103.700 13.990 104.840 14.640 ;
        RECT 105.110 14.570 105.340 16.190 ;
        RECT 106.150 16.180 106.380 16.190 ;
        RECT 106.090 15.620 106.450 16.180 ;
        RECT 105.040 14.010 105.400 14.570 ;
        RECT 103.700 12.840 104.120 13.990 ;
        RECT 104.470 13.970 104.840 13.990 ;
        RECT 104.520 13.950 104.770 13.970 ;
        RECT 105.110 13.940 105.340 14.010 ;
        RECT 106.150 13.940 106.380 15.620 ;
        RECT 107.190 14.540 107.420 16.190 ;
        RECT 107.140 13.980 107.500 14.540 ;
        RECT 107.190 13.940 107.420 13.980 ;
        RECT 108.460 13.800 108.790 16.350 ;
        RECT 111.460 16.340 114.850 16.610 ;
        RECT 117.480 16.340 120.870 16.610 ;
        RECT 111.480 16.330 112.190 16.340 ;
        RECT 112.520 16.330 113.230 16.340 ;
        RECT 110.630 14.530 110.870 14.590 ;
        RECT 105.390 13.530 108.790 13.800 ;
        RECT 109.890 14.500 110.370 14.510 ;
        RECT 110.560 14.500 110.940 14.530 ;
        RECT 111.200 14.520 111.430 16.170 ;
        RECT 112.160 15.730 112.550 16.180 ;
        RECT 109.890 13.950 110.940 14.500 ;
        RECT 111.120 13.970 111.510 14.520 ;
        RECT 109.890 12.840 110.370 13.950 ;
        RECT 110.560 13.940 110.940 13.950 ;
        RECT 110.630 13.910 110.870 13.940 ;
        RECT 111.200 13.920 111.430 13.970 ;
        RECT 112.240 13.920 112.470 15.730 ;
        RECT 113.280 14.460 113.510 16.170 ;
        RECT 113.220 13.960 113.590 14.460 ;
        RECT 113.280 13.920 113.510 13.960 ;
        RECT 114.520 13.780 114.850 16.340 ;
        RECT 116.570 14.480 116.900 14.530 ;
        RECT 117.210 14.500 117.440 16.180 ;
        RECT 118.180 15.730 118.550 16.180 ;
        RECT 115.700 13.930 116.920 14.480 ;
        RECT 117.140 14.000 117.510 14.500 ;
        RECT 117.210 13.930 117.440 14.000 ;
        RECT 118.250 13.930 118.480 15.730 ;
        RECT 119.290 14.490 119.520 16.180 ;
        RECT 119.210 13.990 119.580 14.490 ;
        RECT 119.290 13.930 119.520 13.990 ;
        RECT 111.450 13.510 114.850 13.780 ;
        RECT 115.710 12.860 116.350 13.930 ;
        RECT 116.570 13.910 116.900 13.930 ;
        RECT 120.540 13.790 120.870 16.340 ;
        RECT 117.470 13.520 120.870 13.790 ;
        RECT 122.970 12.860 123.600 12.880 ;
        RECT 115.710 12.840 123.600 12.860 ;
        RECT 103.700 12.510 123.600 12.840 ;
        RECT 115.710 12.500 123.600 12.510 ;
        RECT 120.640 11.920 121.140 11.930 ;
        RECT 105.270 11.490 121.140 11.920 ;
        RECT 104.450 8.950 104.810 9.010 ;
        RECT 105.070 8.960 105.300 11.330 ;
        RECT 106.160 11.310 106.390 11.330 ;
        RECT 106.090 10.790 106.470 11.310 ;
        RECT 104.430 8.110 104.830 8.950 ;
        RECT 104.990 8.120 105.390 8.960 ;
        RECT 104.450 8.050 104.810 8.110 ;
        RECT 105.070 8.080 105.300 8.120 ;
        RECT 106.160 8.080 106.390 10.790 ;
        RECT 107.250 8.970 107.480 11.330 ;
        RECT 110.480 8.970 110.840 9.030 ;
        RECT 111.170 9.000 111.400 11.330 ;
        RECT 112.180 10.780 112.590 11.340 ;
        RECT 107.150 8.130 107.550 8.970 ;
        RECT 110.460 8.130 110.860 8.970 ;
        RECT 111.050 8.160 111.450 9.000 ;
        RECT 107.250 8.080 107.480 8.130 ;
        RECT 110.480 8.070 110.840 8.130 ;
        RECT 111.170 8.080 111.400 8.160 ;
        RECT 112.260 8.080 112.490 10.780 ;
        RECT 113.350 8.940 113.580 11.330 ;
        RECT 113.260 8.100 113.660 8.940 ;
        RECT 116.630 8.820 116.960 8.880 ;
        RECT 117.250 8.820 117.480 11.350 ;
        RECT 118.340 11.260 118.570 11.350 ;
        RECT 118.320 10.690 118.710 11.260 ;
        RECT 116.610 8.170 116.980 8.820 ;
        RECT 117.170 8.170 117.540 8.820 ;
        RECT 116.630 8.110 116.960 8.170 ;
        RECT 117.250 8.100 117.480 8.170 ;
        RECT 118.340 8.100 118.570 10.690 ;
        RECT 119.430 8.760 119.660 11.350 ;
        RECT 120.640 10.700 121.140 11.490 ;
        RECT 125.900 10.700 126.860 18.510 ;
        RECT 140.400 18.080 140.860 18.110 ;
        RECT 141.230 18.080 142.410 18.100 ;
        RECT 140.400 18.070 142.410 18.080 ;
        RECT 143.260 18.070 143.540 18.080 ;
        RECT 138.420 17.620 139.260 17.710 ;
        RECT 140.400 17.680 143.540 18.070 ;
        RECT 140.400 17.670 141.230 17.680 ;
        RECT 140.400 17.620 140.860 17.670 ;
        RECT 142.410 17.660 143.540 17.680 ;
        RECT 138.060 17.560 140.860 17.620 ;
        RECT 138.010 17.490 140.860 17.560 ;
        RECT 138.000 17.240 140.860 17.490 ;
        RECT 141.535 17.420 141.765 17.525 ;
        RECT 138.050 17.225 138.340 17.240 ;
        RECT 138.810 17.200 140.860 17.240 ;
        RECT 137.785 16.940 138.015 17.065 ;
        RECT 137.630 16.370 138.120 16.940 ;
        RECT 137.785 15.065 138.015 16.370 ;
        RECT 138.375 15.760 138.605 17.065 ;
        RECT 138.160 15.270 138.790 15.760 ;
        RECT 139.470 15.380 140.860 17.200 ;
        RECT 141.250 16.680 141.960 17.420 ;
        RECT 141.535 15.525 141.765 16.680 ;
        RECT 142.125 16.280 142.355 17.525 ;
        RECT 143.260 17.260 143.540 17.660 ;
        RECT 141.920 15.730 142.660 16.280 ;
        RECT 143.260 16.090 143.960 17.260 ;
        RECT 148.630 17.130 149.560 17.150 ;
        RECT 148.630 16.870 151.850 17.130 ;
        RECT 148.630 16.750 153.245 16.870 ;
        RECT 147.200 16.700 153.245 16.750 ;
        RECT 143.260 15.950 145.530 16.090 ;
        RECT 143.260 15.750 145.560 15.950 ;
        RECT 142.125 15.525 142.355 15.730 ;
        RECT 139.470 15.340 142.090 15.380 ;
        RECT 143.260 15.340 143.960 15.750 ;
        RECT 145.100 15.720 145.560 15.750 ;
        RECT 147.200 15.760 149.610 16.700 ;
        RECT 151.285 16.640 153.245 16.700 ;
        RECT 151.005 15.960 151.235 16.435 ;
        RECT 144.820 15.480 145.050 15.560 ;
        RECT 138.375 15.065 138.605 15.270 ;
        RECT 139.470 14.970 143.960 15.340 ;
        RECT 144.650 15.010 145.160 15.480 ;
        RECT 145.610 15.370 145.840 15.560 ;
        RECT 139.470 14.960 140.860 14.970 ;
        RECT 139.460 14.940 140.860 14.960 ;
        RECT 138.050 14.890 138.340 14.905 ;
        RECT 139.460 14.900 140.570 14.940 ;
        RECT 142.030 14.930 143.960 14.970 ;
        RECT 139.460 14.890 139.600 14.900 ;
        RECT 143.500 14.890 143.960 14.930 ;
        RECT 138.000 14.660 139.600 14.890 ;
        RECT 138.070 14.580 139.600 14.660 ;
        RECT 143.720 14.690 143.960 14.890 ;
        RECT 144.820 14.860 145.050 15.010 ;
        RECT 145.580 14.900 146.270 15.370 ;
        RECT 147.200 15.350 149.750 15.760 ;
        RECT 150.830 15.560 151.350 15.960 ;
        RECT 153.050 15.570 153.840 16.470 ;
        RECT 155.620 16.440 155.910 16.500 ;
        RECT 155.620 16.400 157.090 16.440 ;
        RECT 154.640 15.680 157.090 16.400 ;
        RECT 151.005 15.435 151.235 15.560 ;
        RECT 153.295 15.435 153.525 15.570 ;
        RECT 148.630 15.280 149.750 15.350 ;
        RECT 148.630 15.230 151.890 15.280 ;
        RECT 148.630 15.000 153.245 15.230 ;
        RECT 154.500 15.160 157.090 15.680 ;
        RECT 155.620 15.110 157.090 15.160 ;
        RECT 155.620 15.040 155.910 15.110 ;
        RECT 145.610 14.860 145.840 14.900 ;
        RECT 148.710 14.880 152.040 15.000 ;
        RECT 148.750 14.860 152.040 14.880 ;
        RECT 145.100 14.690 145.560 14.700 ;
        RECT 143.720 14.470 145.560 14.690 ;
        RECT 151.890 14.670 152.040 14.860 ;
        RECT 141.850 14.040 142.430 14.410 ;
        RECT 143.720 14.350 145.550 14.470 ;
        RECT 141.970 14.030 142.350 14.040 ;
        RECT 146.750 14.010 147.610 14.160 ;
        RECT 154.680 14.010 155.340 14.110 ;
        RECT 137.970 13.040 138.660 13.880 ;
        RECT 141.220 13.830 141.670 13.850 ;
        RECT 142.570 13.830 143.090 13.930 ;
        RECT 141.220 13.580 143.090 13.830 ;
        RECT 141.220 13.490 142.780 13.580 ;
        RECT 141.430 13.050 142.780 13.490 ;
        RECT 143.930 13.150 145.130 13.770 ;
        RECT 146.750 13.550 155.340 14.010 ;
        RECT 141.430 12.940 143.090 13.050 ;
        RECT 141.260 12.690 143.090 12.940 ;
        RECT 145.800 12.710 146.350 13.350 ;
        RECT 147.360 12.890 150.370 13.120 ;
        RECT 147.360 12.780 154.540 12.890 ;
        RECT 141.260 12.650 141.700 12.690 ;
        RECT 142.600 12.630 143.090 12.690 ;
        RECT 147.270 12.680 154.540 12.780 ;
        RECT 147.270 12.530 148.420 12.680 ;
        RECT 149.580 12.660 154.540 12.680 ;
        RECT 147.270 12.510 148.290 12.530 ;
        RECT 147.290 12.280 148.290 12.510 ;
        RECT 154.680 12.500 155.340 13.550 ;
        RECT 146.930 11.670 148.290 12.280 ;
        RECT 149.300 12.270 149.530 12.500 ;
        RECT 149.140 11.830 149.740 12.270 ;
        RECT 146.930 11.340 148.350 11.670 ;
        RECT 149.300 11.500 149.530 11.830 ;
        RECT 154.590 11.620 155.340 12.500 ;
        RECT 154.590 11.500 154.820 11.620 ;
        RECT 146.930 11.110 154.540 11.340 ;
        RECT 146.930 10.920 150.400 11.110 ;
        RECT 147.390 10.900 150.400 10.920 ;
        RECT 120.640 9.750 126.860 10.700 ;
        RECT 119.370 8.110 119.740 8.760 ;
        RECT 119.430 8.100 119.660 8.110 ;
        RECT 113.350 8.080 113.580 8.100 ;
        RECT 117.530 7.930 118.290 7.940 ;
        RECT 118.620 7.930 119.380 7.940 ;
        RECT 120.640 7.930 121.140 9.750 ;
        RECT 105.290 7.540 121.140 7.930 ;
        RECT 105.290 7.500 121.110 7.540 ;
        RECT 109.100 6.060 110.210 6.830 ;
        RECT 109.170 5.920 110.170 6.060 ;
        RECT 109.170 4.790 110.430 5.920 ;
        RECT 109.290 3.470 110.430 4.790 ;
        RECT 108.400 2.630 110.960 3.470 ;
      LAYER met2 ;
        RECT 42.120 223.240 43.620 224.360 ;
        RECT 45.480 223.310 48.340 223.730 ;
        RECT 46.520 222.570 50.740 223.020 ;
        RECT 6.790 221.260 9.810 222.180 ;
        RECT 46.970 221.070 47.270 222.570 ;
        RECT 60.840 220.840 63.250 221.260 ;
        RECT 46.970 217.670 47.270 220.770 ;
        RECT 55.010 218.590 56.140 220.310 ;
        RECT 76.525 219.450 79.210 219.480 ;
        RECT 65.010 218.770 67.680 219.210 ;
        RECT 44.390 215.900 45.790 216.540 ;
        RECT 17.250 214.450 17.710 214.860 ;
        RECT 17.310 213.580 17.630 214.450 ;
        RECT 30.080 214.290 30.510 214.770 ;
        RECT 17.310 213.430 17.640 213.580 ;
        RECT 17.320 213.110 17.640 213.430 ;
        RECT 30.110 213.570 30.470 214.290 ;
        RECT 30.950 214.280 31.620 215.480 ;
        RECT 41.960 214.410 42.430 214.860 ;
        RECT 46.910 214.700 47.380 217.670 ;
        RECT 67.340 216.650 67.680 218.770 ;
        RECT 63.880 216.360 67.680 216.650 ;
        RECT 63.880 215.480 64.220 216.360 ;
        RECT 69.330 216.030 69.660 219.230 ;
        RECT 76.525 218.710 79.610 219.450 ;
        RECT 109.820 218.870 111.200 219.510 ;
        RECT 140.030 219.170 140.630 222.060 ;
        RECT 134.670 218.410 135.130 218.690 ;
        RECT 134.770 218.000 135.080 218.410 ;
        RECT 64.580 215.810 64.920 215.890 ;
        RECT 64.580 215.520 67.680 215.810 ;
        RECT 64.580 215.480 64.920 215.520 ;
        RECT 42.010 213.580 42.360 214.410 ;
        RECT 30.110 213.120 30.460 213.570 ;
        RECT 42.020 213.180 42.360 213.580 ;
        RECT 44.120 214.120 46.410 214.210 ;
        RECT 48.910 214.120 50.610 214.420 ;
        RECT 11.850 212.570 12.110 212.950 ;
        RECT 18.590 212.590 18.870 212.960 ;
        RECT 24.640 212.580 24.920 213.020 ;
        RECT 30.940 212.570 31.220 213.020 ;
        RECT 36.550 212.590 36.900 213.040 ;
        RECT 42.860 212.610 43.180 213.080 ;
        RECT 44.120 212.710 50.610 214.120 ;
        RECT 44.120 212.670 46.410 212.710 ;
        RECT 48.910 212.140 50.610 212.710 ;
        RECT 54.210 211.790 55.610 212.940 ;
        RECT 55.750 212.690 56.100 212.740 ;
        RECT 60.060 212.690 60.450 212.740 ;
        RECT 55.750 212.090 60.450 212.690 ;
        RECT 67.340 212.480 67.680 215.520 ;
        RECT 68.660 215.430 69.660 216.030 ;
        RECT 55.750 212.040 56.100 212.090 ;
        RECT 60.060 212.020 60.450 212.090 ;
        RECT 65.210 212.060 67.680 212.480 ;
        RECT 69.330 212.190 69.660 215.430 ;
        RECT 77.670 213.710 78.380 217.700 ;
        RECT 128.460 216.250 129.220 217.110 ;
        RECT 132.460 217.030 132.970 217.070 ;
        RECT 132.460 217.020 133.840 217.030 ;
        RECT 132.460 216.490 134.190 217.020 ;
        RECT 132.460 216.470 133.840 216.490 ;
        RECT 132.460 216.410 132.970 216.470 ;
        RECT 134.760 216.280 135.090 218.000 ;
        RECT 134.730 215.890 135.150 216.280 ;
        RECT 76.390 211.880 79.560 212.630 ;
        RECT 106.500 212.270 107.790 213.660 ;
        RECT 81.410 209.910 85.680 210.050 ;
        RECT 8.110 209.610 85.680 209.910 ;
        RECT 8.110 202.840 8.410 209.610 ;
        RECT 81.410 209.520 85.680 209.610 ;
        RECT 9.120 206.510 12.210 209.110 ;
        RECT 19.270 206.830 25.300 208.840 ;
        RECT 75.300 206.630 78.390 209.160 ;
        RECT 82.170 206.610 83.990 209.050 ;
        RECT 84.610 203.680 85.230 206.260 ;
        RECT 115.040 205.620 117.310 209.190 ;
        RECT 129.850 206.140 130.950 208.270 ;
        RECT 134.630 208.250 135.090 208.530 ;
        RECT 132.430 206.880 132.940 206.990 ;
        RECT 133.750 206.880 134.160 206.910 ;
        RECT 132.430 206.410 134.160 206.880 ;
        RECT 132.430 206.330 132.940 206.410 ;
        RECT 133.750 206.380 134.160 206.410 ;
        RECT 134.720 205.960 135.010 208.250 ;
        RECT 134.670 205.570 135.090 205.960 ;
        RECT 117.050 203.580 118.380 204.750 ;
        RECT 30.830 203.380 31.170 203.410 ;
        RECT 18.430 203.270 18.790 203.310 ;
        RECT 8.050 199.750 8.860 202.840 ;
        RECT 18.420 199.990 18.800 203.270 ;
        RECT 30.810 200.400 31.170 203.380 ;
        RECT 43.090 202.810 43.720 203.340 ;
        RECT 30.810 200.030 31.230 200.400 ;
        RECT 43.150 200.070 43.720 202.810 ;
        RECT 43.160 200.010 43.610 200.070 ;
        RECT 55.580 199.510 58.080 202.110 ;
        RECT 85.410 199.490 87.170 202.130 ;
        RECT 49.100 196.550 50.300 199.010 ;
        RECT 134.640 198.140 135.100 198.420 ;
        RECT 134.700 198.080 135.100 198.140 ;
        RECT 132.810 196.840 133.890 196.850 ;
        RECT 132.390 196.800 133.890 196.840 ;
        RECT 132.390 196.270 134.230 196.800 ;
        RECT 134.760 196.750 135.100 198.080 ;
        RECT 134.700 196.350 135.140 196.750 ;
        RECT 134.700 196.340 135.090 196.350 ;
        RECT 132.390 196.200 133.890 196.270 ;
        RECT 132.390 196.180 132.900 196.200 ;
        RECT 134.760 195.860 135.090 196.340 ;
        RECT 134.760 195.810 135.140 195.860 ;
        RECT 134.760 195.770 135.190 195.810 ;
        RECT 94.330 194.460 95.330 195.560 ;
        RECT 97.750 193.280 98.380 195.010 ;
        RECT 97.740 192.850 98.380 193.280 ;
        RECT 103.620 193.190 104.330 194.740 ;
        RECT 110.760 194.370 111.630 195.590 ;
        RECT 134.770 195.420 135.190 195.770 ;
        RECT 103.610 193.160 104.330 193.190 ;
        RECT 103.610 192.640 104.300 193.160 ;
        RECT 105.250 192.340 105.690 192.390 ;
        RECT 108.700 192.340 109.140 192.370 ;
        RECT 105.250 191.860 109.140 192.340 ;
        RECT 105.250 191.830 105.690 191.860 ;
        RECT 108.700 191.810 109.140 191.860 ;
        RECT 99.740 189.870 100.120 190.190 ;
        RECT 99.740 188.700 100.130 189.870 ;
        RECT 136.330 189.630 138.020 193.530 ;
        RECT 97.160 188.370 100.130 188.700 ;
        RECT 93.420 185.580 94.420 186.680 ;
        RECT 97.170 186.520 97.530 188.370 ;
        RECT 94.640 186.460 95.080 186.510 ;
        RECT 97.090 186.480 97.530 186.520 ;
        RECT 95.960 186.460 97.530 186.480 ;
        RECT 94.640 185.820 97.530 186.460 ;
        RECT 94.640 185.780 95.080 185.820 ;
        RECT 95.960 185.810 97.530 185.820 ;
        RECT 97.090 185.790 97.530 185.810 ;
        RECT 103.570 188.320 104.260 188.820 ;
        RECT 103.570 185.770 104.310 188.320 ;
        RECT 125.230 187.780 129.570 188.970 ;
        RECT 103.580 185.660 104.310 185.770 ;
        RECT 110.690 185.750 111.610 186.860 ;
        RECT 103.660 185.620 104.240 185.660 ;
        RECT 48.890 183.330 50.690 185.190 ;
        RECT 48.850 176.950 52.440 181.650 ;
        RECT 132.650 178.110 137.990 180.650 ;
        RECT 143.770 175.070 144.170 178.490 ;
        RECT 147.450 175.020 147.970 178.630 ;
        RECT 40.590 153.870 47.630 155.370 ;
        RECT 1.010 148.870 11.810 153.540 ;
        RECT 72.500 150.340 82.530 151.380 ;
        RECT 101.860 150.540 103.120 151.950 ;
        RECT 85.110 150.340 86.500 150.410 ;
        RECT 72.500 150.310 86.500 150.340 ;
        RECT 72.500 150.260 86.510 150.310 ;
        RECT 72.670 149.830 86.510 150.260 ;
        RECT 72.750 149.610 75.740 149.830 ;
        RECT 85.110 149.810 86.500 149.830 ;
        RECT 84.000 149.630 84.380 149.680 ;
        RECT 51.780 147.090 55.790 149.380 ;
        RECT 83.980 149.190 84.380 149.630 ;
        RECT 77.120 148.650 77.590 148.690 ;
        RECT 77.110 148.590 78.110 148.650 ;
        RECT 83.980 148.590 84.370 149.190 ;
        RECT 77.110 148.190 84.370 148.590 ;
        RECT 62.855 148.110 63.315 148.160 ;
        RECT 62.845 147.730 63.315 148.110 ;
        RECT 59.230 146.930 59.940 146.940 ;
        RECT 62.845 146.930 63.305 147.730 ;
        RECT 77.110 147.590 78.110 148.190 ;
        RECT 77.120 147.540 77.590 147.590 ;
        RECT 69.250 147.400 70.520 147.470 ;
        RECT 72.770 147.400 73.970 147.460 ;
        RECT 56.360 145.760 57.500 146.600 ;
        RECT 59.230 146.590 63.310 146.930 ;
        RECT 69.250 146.900 73.970 147.400 ;
        RECT 81.130 147.430 81.390 147.490 ;
        RECT 81.130 147.050 81.710 147.430 ;
        RECT 59.230 145.180 59.940 146.590 ;
        RECT 60.290 145.850 61.280 146.440 ;
        RECT 69.250 146.080 70.520 146.900 ;
        RECT 72.770 146.880 73.970 146.900 ;
        RECT 59.220 145.020 59.940 145.180 ;
        RECT 59.220 144.250 59.960 145.020 ;
        RECT 66.360 144.800 66.700 144.860 ;
        RECT 59.220 143.080 59.900 144.250 ;
        RECT 66.330 143.310 66.710 144.800 ;
        RECT 77.140 144.700 78.110 144.790 ;
        RECT 77.140 144.090 78.140 144.700 ;
        RECT 81.440 144.490 81.710 147.050 ;
        RECT 85.150 144.860 86.700 147.420 ;
        RECT 88.730 146.870 89.570 147.970 ;
        RECT 90.790 147.030 91.580 147.890 ;
        RECT 81.440 144.420 81.700 144.490 ;
        RECT 77.140 143.740 84.900 144.090 ;
        RECT 77.140 143.670 78.140 143.740 ;
        RECT 70.890 143.380 71.260 143.480 ;
        RECT 70.730 143.310 71.260 143.380 ;
        RECT 66.330 143.180 71.260 143.310 ;
        RECT 59.210 142.750 63.710 143.080 ;
        RECT 66.330 142.810 71.370 143.180 ;
        RECT 77.120 143.080 78.140 143.670 ;
        RECT 84.530 143.290 84.900 143.740 ;
        RECT 66.330 142.790 68.940 142.810 ;
        RECT 63.270 140.740 63.710 142.750 ;
        RECT 68.540 141.460 68.940 142.790 ;
        RECT 70.730 142.710 71.260 142.810 ;
        RECT 70.890 142.630 71.260 142.710 ;
        RECT 77.120 142.590 78.120 143.080 ;
        RECT 68.510 140.740 68.970 141.460 ;
        RECT 88.310 141.040 88.620 141.970 ;
        RECT 63.260 140.370 63.710 140.740 ;
        RECT 88.850 140.610 89.570 146.870 ;
        RECT 90.800 142.720 91.580 147.030 ;
        RECT 98.230 145.560 99.410 145.620 ;
        RECT 96.900 145.010 99.410 145.560 ;
        RECT 90.230 142.240 91.820 142.720 ;
        RECT 88.850 140.580 90.250 140.610 ;
        RECT 88.850 138.540 90.260 140.580 ;
        RECT 91.250 139.120 92.320 140.620 ;
        RECT 88.850 137.990 92.150 138.540 ;
        RECT 79.440 136.950 79.730 137.100 ;
        RECT 70.090 136.490 70.360 136.590 ;
        RECT 73.890 136.490 74.200 136.550 ;
        RECT 70.090 136.250 74.200 136.490 ;
        RECT 70.090 136.170 70.360 136.250 ;
        RECT 73.890 136.150 74.200 136.250 ;
        RECT 79.430 135.490 79.730 136.950 ;
        RECT 82.250 136.420 83.810 137.580 ;
        RECT 94.050 137.070 94.870 137.580 ;
        RECT 96.910 137.070 97.470 145.010 ;
        RECT 98.230 144.970 99.410 145.010 ;
        RECT 98.400 141.060 99.340 141.610 ;
        RECT 97.840 138.590 99.310 139.290 ;
        RECT 94.050 136.720 97.470 137.070 ;
        RECT 79.430 135.240 81.030 135.490 ;
        RECT 80.720 133.650 81.030 135.240 ;
        RECT 82.250 135.050 89.350 136.420 ;
        RECT 94.050 136.230 94.870 136.720 ;
        RECT 96.910 136.700 97.470 136.720 ;
        RECT 82.250 134.800 83.810 135.050 ;
        RECT 79.400 133.190 79.720 133.550 ;
        RECT 80.720 133.190 81.040 133.650 ;
        RECT 70.010 132.960 70.290 133.060 ;
        RECT 70.010 132.950 70.780 132.960 ;
        RECT 73.850 132.950 74.140 133.010 ;
        RECT 70.010 132.670 74.140 132.950 ;
        RECT 70.010 132.580 70.290 132.670 ;
        RECT 73.850 132.620 74.140 132.670 ;
        RECT 79.410 131.970 79.700 133.190 ;
        RECT 111.630 131.970 114.370 134.600 ;
        RECT 79.410 131.770 81.010 131.970 ;
        RECT 80.790 130.130 81.010 131.770 ;
        RECT 80.740 129.690 81.080 130.130 ;
        RECT 69.930 129.480 70.250 129.530 ;
        RECT 69.920 129.160 74.240 129.480 ;
        RECT 69.930 129.110 70.250 129.160 ;
        RECT 73.920 129.110 74.240 129.160 ;
        RECT 81.410 128.510 83.550 131.140 ;
        RECT 85.220 129.720 87.570 131.320 ;
        RECT 108.770 129.730 111.040 131.370 ;
        RECT 1.010 32.995 5.080 33.890 ;
        RECT 113.100 32.995 118.190 33.200 ;
        RECT 1.010 32.980 142.075 32.995 ;
        RECT 1.010 31.725 142.130 32.980 ;
        RECT 1.010 30.360 5.080 31.725 ;
        RECT 113.100 31.650 118.190 31.725 ;
        RECT 100.630 29.460 101.350 29.480 ;
        RECT 100.630 29.430 115.740 29.460 ;
        RECT 100.630 29.060 115.830 29.430 ;
        RECT 140.180 29.300 142.130 31.725 ;
        RECT 143.740 30.320 144.230 32.790 ;
        RECT 147.350 30.260 148.010 32.770 ;
        RECT 144.130 29.300 145.850 29.960 ;
        RECT 152.020 29.330 152.820 29.460 ;
        RECT 147.550 29.300 152.820 29.330 ;
        RECT 100.630 28.700 115.840 29.060 ;
        RECT 100.630 20.920 101.350 28.700 ;
        RECT 103.680 22.760 104.140 28.700 ;
        RECT 106.220 27.510 106.510 27.560 ;
        RECT 109.010 27.510 109.270 27.520 ;
        RECT 111.850 27.510 112.140 27.530 ;
        RECT 115.080 27.510 115.840 28.700 ;
        RECT 140.180 28.060 152.820 29.300 ;
        RECT 140.550 28.040 152.770 28.060 ;
        RECT 116.400 27.510 116.700 27.550 ;
        RECT 117.000 27.510 117.260 27.530 ;
        RECT 121.530 27.510 121.840 27.580 ;
        RECT 122.140 27.510 122.400 27.560 ;
        RECT 124.330 27.510 124.590 27.560 ;
        RECT 106.220 26.880 124.680 27.510 ;
        RECT 106.220 26.810 106.510 26.880 ;
        RECT 106.790 26.770 107.050 26.880 ;
        RECT 109.010 26.790 109.270 26.880 ;
        RECT 111.320 26.650 111.610 26.880 ;
        RECT 111.850 26.730 112.140 26.880 ;
        RECT 114.110 26.690 114.400 26.880 ;
        RECT 116.400 26.660 116.700 26.880 ;
        RECT 117.000 26.800 117.260 26.880 ;
        RECT 119.190 26.760 119.450 26.880 ;
        RECT 121.530 26.710 121.840 26.880 ;
        RECT 122.140 26.830 122.400 26.880 ;
        RECT 124.330 26.830 124.590 26.880 ;
        RECT 140.550 26.570 141.760 28.040 ;
        RECT 143.470 27.870 145.130 28.040 ;
        RECT 140.390 26.370 141.760 26.570 ;
        RECT 140.080 26.270 141.760 26.370 ;
        RECT 118.080 25.100 118.380 25.120 ;
        RECT 112.970 24.970 113.250 24.990 ;
        RECT 107.850 24.350 108.140 24.920 ;
        RECT 107.850 24.270 108.150 24.350 ;
        RECT 103.720 22.710 104.140 22.760 ;
        RECT 100.630 20.910 101.650 20.920 ;
        RECT 99.300 20.870 99.620 20.910 ;
        RECT 100.380 20.870 101.650 20.910 ;
        RECT 99.290 20.440 101.710 20.870 ;
        RECT 99.300 20.380 99.620 20.440 ;
        RECT 100.380 20.380 100.700 20.440 ;
        RECT 101.330 20.390 101.650 20.440 ;
        RECT 103.720 20.390 104.110 22.710 ;
        RECT 107.860 22.680 108.150 24.270 ;
        RECT 109.710 22.700 110.140 23.120 ;
        RECT 106.680 22.390 108.150 22.680 ;
        RECT 105.320 20.830 105.640 20.870 ;
        RECT 105.320 20.810 105.650 20.830 ;
        RECT 106.680 20.810 107.040 22.390 ;
        RECT 107.860 22.380 108.150 22.390 ;
        RECT 107.420 20.810 107.740 20.840 ;
        RECT 103.740 20.320 104.000 20.390 ;
        RECT 105.320 20.370 107.780 20.810 ;
        RECT 105.320 20.340 105.640 20.370 ;
        RECT 107.420 20.310 107.740 20.370 ;
        RECT 109.740 20.330 110.130 22.700 ;
        RECT 111.420 20.820 111.690 20.860 ;
        RECT 112.940 20.820 113.310 24.970 ;
        RECT 118.080 24.230 118.490 25.100 ;
        RECT 139.910 25.080 141.760 26.270 ;
        RECT 145.890 26.180 146.760 28.040 ;
        RECT 147.550 28.030 152.770 28.040 ;
        RECT 151.750 27.310 152.770 28.030 ;
        RECT 151.750 27.300 152.780 27.310 ;
        RECT 145.840 25.670 146.760 26.180 ;
        RECT 151.780 26.430 152.780 27.300 ;
        RECT 145.840 25.470 146.280 25.670 ;
        RECT 151.780 25.320 152.820 26.430 ;
        RECT 152.160 25.270 152.500 25.320 ;
        RECT 140.080 25.020 141.760 25.080 ;
        RECT 123.210 24.970 123.500 25.020 ;
        RECT 140.080 24.990 140.670 25.020 ;
        RECT 140.410 24.970 140.670 24.990 ;
        RECT 141.240 24.980 141.640 25.020 ;
        RECT 115.790 22.690 116.220 23.110 ;
        RECT 113.490 20.820 113.760 20.850 ;
        RECT 111.420 20.370 113.760 20.820 ;
        RECT 111.420 20.350 111.690 20.370 ;
        RECT 113.490 20.340 113.760 20.370 ;
        RECT 115.800 20.200 116.190 22.690 ;
        RECT 117.490 20.730 117.750 20.840 ;
        RECT 118.100 20.730 118.490 24.230 ;
        RECT 123.170 20.900 123.500 24.970 ;
        RECT 136.840 22.960 138.210 24.530 ;
        RECT 139.450 22.340 139.930 22.450 ;
        RECT 140.670 22.340 141.150 22.420 ;
        RECT 139.450 21.010 141.220 22.340 ;
        RECT 139.050 20.940 141.220 21.010 ;
        RECT 151.600 21.320 151.970 21.470 ;
        RECT 152.750 21.320 153.120 21.450 ;
        RECT 123.190 20.850 123.450 20.900 ;
        RECT 119.550 20.730 119.810 20.810 ;
        RECT 117.490 20.210 119.840 20.730 ;
        RECT 117.490 20.200 117.750 20.210 ;
        RECT 115.850 20.180 116.110 20.200 ;
        RECT 119.550 20.170 119.810 20.210 ;
        RECT 99.920 19.360 100.180 19.420 ;
        RECT 100.890 19.360 101.150 19.390 ;
        RECT 99.880 18.930 101.160 19.360 ;
        RECT 104.270 19.250 104.570 19.280 ;
        RECT 106.390 19.250 106.690 19.310 ;
        RECT 99.920 18.900 100.180 18.930 ;
        RECT 100.730 18.870 101.150 18.930 ;
        RECT 96.630 17.010 98.880 18.200 ;
        RECT 100.730 17.880 101.090 18.870 ;
        RECT 104.270 18.850 106.690 19.250 ;
        RECT 104.270 18.740 104.570 18.850 ;
        RECT 106.090 18.770 106.690 18.850 ;
        RECT 110.360 19.290 110.640 19.340 ;
        RECT 116.420 19.310 116.680 19.360 ;
        RECT 118.500 19.310 118.760 19.360 ;
        RECT 112.440 19.290 112.720 19.300 ;
        RECT 110.360 18.780 112.730 19.290 ;
        RECT 116.420 18.800 118.790 19.310 ;
        RECT 121.510 19.020 121.790 19.140 ;
        RECT 122.030 19.020 122.380 19.110 ;
        RECT 124.220 19.020 124.570 19.050 ;
        RECT 100.720 17.300 101.120 17.880 ;
        RECT 102.200 17.670 102.530 17.730 ;
        RECT 106.090 17.670 106.440 18.770 ;
        RECT 102.200 17.310 106.440 17.670 ;
        RECT 112.200 18.740 112.720 18.780 ;
        RECT 116.420 18.760 116.680 18.800 ;
        RECT 118.180 18.760 118.760 18.800 ;
        RECT 112.200 17.660 112.500 18.740 ;
        RECT 114.530 17.660 114.870 17.710 ;
        RECT 118.180 17.660 118.500 18.760 ;
        RECT 121.500 18.310 124.600 19.020 ;
        RECT 126.870 18.460 128.430 20.290 ;
        RECT 139.050 18.780 140.040 20.940 ;
        RECT 140.670 20.840 141.150 20.940 ;
        RECT 151.600 20.740 153.240 21.320 ;
        RECT 151.600 20.390 153.680 20.740 ;
        RECT 151.600 20.320 151.970 20.390 ;
        RECT 136.940 18.560 140.040 18.780 ;
        RECT 121.510 18.270 121.790 18.310 ;
        RECT 122.030 18.300 122.380 18.310 ;
        RECT 100.730 15.540 101.090 17.300 ;
        RECT 102.200 17.250 102.530 17.310 ;
        RECT 106.090 17.300 106.440 17.310 ;
        RECT 106.100 15.620 106.430 17.300 ;
        RECT 112.190 17.280 112.510 17.660 ;
        RECT 114.520 17.360 118.530 17.660 ;
        RECT 114.530 17.310 114.870 17.360 ;
        RECT 112.200 15.710 112.500 17.280 ;
        RECT 118.180 15.730 118.500 17.360 ;
        RECT 112.210 15.680 112.500 15.710 ;
        RECT 118.230 15.680 118.500 15.730 ;
        RECT 106.140 15.570 106.400 15.620 ;
        RECT 100.790 15.490 101.050 15.540 ;
        RECT 99.730 14.430 100.000 14.490 ;
        RECT 100.280 14.430 100.550 14.460 ;
        RECT 101.240 14.430 101.510 14.470 ;
        RECT 99.700 13.890 101.530 14.430 ;
        RECT 104.520 13.920 104.790 14.690 ;
        RECT 105.090 14.590 105.350 14.620 ;
        RECT 105.090 13.970 107.460 14.590 ;
        RECT 105.090 13.960 105.350 13.970 ;
        RECT 99.730 13.870 100.000 13.890 ;
        RECT 100.280 13.840 100.550 13.890 ;
        RECT 100.750 13.850 101.510 13.890 ;
        RECT 48.970 5.130 52.940 7.460 ;
        RECT 100.750 6.790 101.320 13.850 ;
        RECT 106.120 10.790 106.420 13.970 ;
        RECT 107.190 13.930 107.450 13.970 ;
        RECT 110.610 13.890 110.890 14.580 ;
        RECT 111.170 14.500 111.460 14.570 ;
        RECT 113.270 14.500 113.540 14.510 ;
        RECT 111.170 13.960 113.550 14.500 ;
        RECT 116.600 14.490 116.870 14.520 ;
        RECT 116.540 13.990 116.870 14.490 ;
        RECT 111.170 13.920 111.460 13.960 ;
        RECT 106.140 10.740 106.420 10.790 ;
        RECT 112.210 10.780 112.540 13.960 ;
        RECT 113.270 13.910 113.540 13.960 ;
        RECT 116.600 13.920 116.870 13.990 ;
        RECT 117.190 14.490 117.460 14.550 ;
        RECT 119.260 14.490 119.530 14.540 ;
        RECT 117.190 13.990 119.590 14.490 ;
        RECT 117.190 13.950 117.460 13.990 ;
        RECT 118.350 11.230 118.680 13.990 ;
        RECT 119.260 13.940 119.530 13.990 ;
        RECT 112.230 10.730 112.540 10.780 ;
        RECT 118.370 10.670 118.680 11.230 ;
        RECT 118.370 10.640 118.660 10.670 ;
        RECT 104.480 8.940 104.780 9.000 ;
        RECT 105.040 8.940 105.340 9.010 ;
        RECT 107.200 8.940 107.500 9.020 ;
        RECT 110.510 8.940 110.810 9.020 ;
        RECT 111.100 8.940 111.400 9.050 ;
        RECT 113.310 8.940 113.610 8.990 ;
        RECT 104.420 8.100 119.740 8.940 ;
        RECT 104.480 8.060 104.780 8.100 ;
        RECT 105.040 8.070 105.340 8.100 ;
        RECT 107.200 8.080 107.500 8.100 ;
        RECT 109.140 6.880 110.150 8.100 ;
        RECT 110.510 8.080 110.810 8.100 ;
        RECT 113.310 8.050 113.610 8.100 ;
        RECT 119.420 8.060 119.690 8.100 ;
        RECT 109.140 6.820 110.160 6.880 ;
        RECT 123.010 6.820 123.690 18.310 ;
        RECT 124.220 18.240 124.570 18.310 ;
        RECT 136.930 18.260 140.040 18.560 ;
        RECT 140.860 19.340 142.110 19.360 ;
        RECT 140.860 18.510 142.300 19.340 ;
        RECT 152.500 18.830 153.680 20.390 ;
        RECT 136.930 18.240 139.100 18.260 ;
        RECT 136.930 17.600 137.890 18.240 ;
        RECT 138.060 18.210 139.100 18.240 ;
        RECT 138.520 17.760 139.100 18.210 ;
        RECT 140.860 18.160 142.130 18.510 ;
        RECT 140.860 18.130 141.760 18.160 ;
        RECT 136.930 17.210 137.870 17.600 ;
        RECT 138.470 17.390 139.210 17.760 ;
        RECT 140.860 17.640 141.750 18.130 ;
        RECT 152.520 17.970 153.670 18.830 ;
        RECT 140.860 17.470 141.760 17.640 ;
        RECT 136.930 17.080 137.910 17.210 ;
        RECT 136.930 16.990 138.050 17.080 ;
        RECT 136.930 16.460 138.070 16.990 ;
        RECT 140.860 16.670 141.910 17.470 ;
        RECT 152.520 17.060 153.690 17.970 ;
        RECT 144.800 16.680 145.290 16.690 ;
        RECT 146.360 16.680 147.030 16.710 ;
        RECT 141.300 16.630 141.910 16.670 ;
        RECT 137.410 16.420 138.070 16.460 ;
        RECT 137.680 16.320 138.070 16.420 ;
        RECT 141.970 16.070 142.610 16.330 ;
        RECT 144.780 16.250 147.030 16.680 ;
        RECT 138.190 15.680 138.740 15.810 ;
        RECT 141.970 15.680 142.840 16.070 ;
        RECT 138.190 15.390 139.070 15.680 ;
        RECT 138.190 15.220 139.050 15.390 ;
        RECT 138.340 13.880 139.050 15.220 ;
        RECT 142.110 14.440 142.840 15.680 ;
        RECT 144.800 15.530 145.290 16.250 ;
        RECT 144.700 15.430 145.290 15.530 ;
        RECT 144.700 15.110 145.310 15.430 ;
        RECT 144.700 14.960 145.110 15.110 ;
        RECT 145.630 14.850 146.220 15.420 ;
        RECT 145.630 14.610 146.150 14.850 ;
        RECT 142.020 14.430 142.840 14.440 ;
        RECT 142.020 13.980 142.940 14.430 ;
        RECT 109.140 6.790 123.690 6.820 ;
        RECT 100.750 6.510 123.690 6.790 ;
        RECT 100.780 6.140 123.690 6.510 ;
        RECT 109.150 6.010 123.690 6.140 ;
        RECT 109.430 5.960 123.690 6.010 ;
        RECT 137.940 13.740 139.050 13.880 ;
        RECT 141.270 13.830 141.620 13.900 ;
        RECT 142.110 13.830 143.040 13.980 ;
        RECT 141.270 13.770 143.040 13.830 ;
        RECT 141.270 13.760 143.690 13.770 ;
        RECT 141.270 13.740 143.750 13.760 ;
        RECT 137.940 13.520 143.750 13.740 ;
        RECT 144.200 13.520 144.950 13.720 ;
        RECT 145.600 13.520 146.170 14.610 ;
        RECT 146.360 14.210 147.030 16.250 ;
        RECT 147.260 15.370 148.300 16.630 ;
        RECT 152.490 16.520 153.670 17.060 ;
        RECT 150.880 15.880 151.300 16.010 ;
        RECT 150.880 15.510 151.560 15.880 ;
        RECT 152.490 15.650 153.790 16.520 ;
        RECT 153.100 15.520 153.790 15.650 ;
        RECT 154.550 15.610 155.620 15.730 ;
        RECT 150.980 14.700 151.560 15.510 ;
        RECT 154.520 15.110 155.620 15.610 ;
        RECT 150.980 14.560 151.630 14.700 ;
        RECT 154.520 14.560 155.450 15.110 ;
        RECT 155.830 15.060 157.040 16.490 ;
        RECT 146.360 13.580 147.560 14.210 ;
        RECT 149.220 13.960 155.460 14.560 ;
        RECT 137.940 13.300 146.140 13.520 ;
        RECT 146.800 13.500 147.560 13.580 ;
        RECT 149.260 13.540 155.460 13.960 ;
        RECT 137.940 12.980 146.210 13.300 ;
        RECT 51.660 3.390 52.420 5.130 ;
        RECT 108.450 3.390 110.910 3.520 ;
        RECT 137.940 3.390 138.700 12.980 ;
        RECT 141.270 12.880 146.210 12.980 ;
        RECT 141.270 12.690 143.040 12.880 ;
        RECT 143.600 12.850 143.960 12.880 ;
        RECT 145.930 12.730 146.210 12.880 ;
        RECT 141.270 12.660 141.650 12.690 ;
        RECT 141.310 12.600 141.650 12.660 ;
        RECT 142.650 12.580 143.040 12.690 ;
        RECT 146.980 10.870 148.040 12.330 ;
        RECT 149.270 12.320 150.060 13.540 ;
        RECT 149.190 11.890 150.060 12.320 ;
        RECT 149.190 11.780 149.690 11.890 ;
        RECT 51.660 2.630 138.720 3.390 ;
        RECT 108.450 2.580 110.910 2.630 ;
      LAYER met3 ;
        RECT 68.180 224.370 70.570 224.620 ;
        RECT 42.060 224.120 70.570 224.370 ;
        RECT 83.100 224.280 83.420 224.320 ;
        RECT 42.060 224.070 70.550 224.120 ;
        RECT 42.070 223.265 43.670 224.070 ;
        RECT 83.100 223.980 130.160 224.280 ;
        RECT 83.100 223.940 83.420 223.980 ;
        RECT 71.610 223.760 74.290 223.920 ;
        RECT 45.380 223.460 74.290 223.760 ;
        RECT 45.430 223.335 48.390 223.460 ;
        RECT 79.370 223.450 79.690 223.490 ;
        RECT 128.140 223.450 128.810 223.460 ;
        RECT 50.740 223.060 67.420 223.160 ;
        RECT 79.370 223.150 128.810 223.450 ;
        RECT 129.460 223.330 130.160 223.980 ;
        RECT 79.370 223.110 79.690 223.150 ;
        RECT 50.460 222.995 67.420 223.060 ;
        RECT 3.950 222.590 4.330 222.910 ;
        RECT 46.470 222.860 67.420 222.995 ;
        RECT 46.470 222.595 51.450 222.860 ;
        RECT 65.130 222.840 67.420 222.860 ;
        RECT 3.990 218.510 4.290 222.590 ;
        RECT 50.460 222.560 51.450 222.595 ;
        RECT 60.700 222.510 62.050 222.530 ;
        RECT 64.170 222.510 65.750 222.530 ;
        RECT 60.700 222.210 65.750 222.510 ;
        RECT 128.140 222.390 128.810 223.150 ;
        RECT 64.170 222.190 65.750 222.210 ;
        RECT 6.740 222.060 9.860 222.155 ;
        RECT 6.660 221.850 9.860 222.060 ;
        RECT 136.110 221.850 136.890 222.130 ;
        RECT 6.660 221.760 136.890 221.850 ;
        RECT 6.740 221.550 136.890 221.760 ;
        RECT 6.740 221.285 9.860 221.550 ;
        RECT 136.110 221.530 136.890 221.550 ;
        RECT 16.800 220.470 17.120 220.510 ;
        RECT 26.000 220.470 26.460 221.220 ;
        RECT 40.520 220.770 54.490 221.070 ;
        RECT 60.790 220.865 63.300 221.235 ;
        RECT 40.520 220.710 42.450 220.770 ;
        RECT 16.800 220.170 26.460 220.470 ;
        RECT 16.800 220.130 17.120 220.170 ;
        RECT 26.000 220.100 26.460 220.170 ;
        RECT 54.110 219.880 54.540 220.770 ;
        RECT 22.350 219.130 22.730 219.140 ;
        RECT 48.950 219.130 50.580 219.360 ;
        RECT 22.350 218.830 50.580 219.130 ;
        RECT 22.350 218.820 22.730 218.830 ;
        RECT 48.950 218.510 50.580 218.830 ;
        RECT 54.960 218.615 56.190 220.285 ;
        RECT 109.770 218.895 111.250 219.485 ;
        RECT 139.980 219.195 140.680 222.035 ;
        RECT 3.990 218.210 50.580 218.510 ;
        RECT 48.950 218.120 50.580 218.210 ;
        RECT 44.340 216.250 45.840 216.515 ;
        RECT 31.130 215.950 45.840 216.250 ;
        RECT 31.130 215.455 31.430 215.950 ;
        RECT 44.340 215.925 45.840 215.950 ;
        RECT 30.900 214.305 31.670 215.455 ;
        RECT 48.730 212.050 50.920 214.530 ;
        RECT 77.620 213.735 78.430 217.675 ;
        RECT 128.410 216.275 129.270 217.085 ;
        RECT 77.710 213.530 78.370 213.735 ;
        RECT 54.160 211.815 55.660 212.915 ;
        RECT 106.530 212.345 107.720 213.525 ;
        RECT 95.830 211.810 96.580 211.920 ;
        RECT 119.550 211.810 120.380 211.990 ;
        RECT 78.820 211.685 79.520 211.760 ;
        RECT 88.560 211.685 89.040 211.760 ;
        RECT 78.820 211.385 89.040 211.685 ;
        RECT 78.820 211.300 79.520 211.385 ;
        RECT 88.560 211.320 89.040 211.385 ;
        RECT 95.830 211.510 120.380 211.810 ;
        RECT 79.740 210.960 80.180 211.050 ;
        RECT 84.860 210.960 85.300 210.980 ;
        RECT 79.740 210.660 85.300 210.960 ;
        RECT 79.740 210.570 80.180 210.660 ;
        RECT 84.860 210.500 85.300 210.660 ;
        RECT 92.140 210.960 93.090 211.300 ;
        RECT 95.830 211.270 96.580 211.510 ;
        RECT 119.550 211.270 120.380 211.510 ;
        RECT 92.140 210.810 93.240 210.960 ;
        RECT 120.890 210.810 122.050 210.830 ;
        RECT 92.140 210.510 122.050 210.810 ;
        RECT 92.140 210.280 93.090 210.510 ;
        RECT 120.890 210.310 122.050 210.510 ;
        RECT 81.360 209.910 85.730 210.025 ;
        RECT 130.950 209.910 131.760 211.380 ;
        RECT 81.360 209.610 131.770 209.910 ;
        RECT 81.360 209.545 85.730 209.610 ;
        RECT 8.990 206.440 12.450 209.190 ;
        RECT 42.665 209.120 45.155 209.135 ;
        RECT 48.990 209.120 50.510 209.160 ;
        RECT 75.250 209.120 78.440 209.135 ;
        RECT 114.990 209.120 117.360 209.165 ;
        RECT 19.220 206.855 25.350 208.815 ;
        RECT 42.620 206.620 117.360 209.120 ;
        RECT 42.660 206.610 45.740 206.620 ;
        RECT 42.665 206.585 45.155 206.610 ;
        RECT 48.990 206.570 50.510 206.620 ;
        RECT 84.560 203.705 85.280 206.235 ;
        RECT 114.990 205.645 117.360 206.620 ;
        RECT 129.800 206.165 131.000 208.245 ;
        RECT 117.000 203.605 118.430 204.725 ;
        RECT 48.930 202.060 52.620 202.090 ;
        RECT 55.530 202.060 58.130 202.085 ;
        RECT 85.360 202.060 87.220 202.105 ;
        RECT 48.930 199.560 87.360 202.060 ;
        RECT 55.530 199.535 58.130 199.560 ;
        RECT 85.360 199.515 87.220 199.560 ;
        RECT 49.050 196.575 50.350 198.985 ;
        RECT 79.700 193.680 80.270 196.770 ;
        RECT 94.280 194.485 95.380 195.535 ;
        RECT 110.710 194.395 111.680 195.565 ;
        RECT 79.730 193.670 80.250 193.680 ;
        RECT 136.410 193.505 138.040 193.520 ;
        RECT 136.280 189.655 138.070 193.505 ;
        RECT 136.280 189.480 138.040 189.655 ;
        RECT 125.090 188.990 128.090 189.170 ;
        RECT 125.090 188.945 128.200 188.990 ;
        RECT 125.090 187.805 129.620 188.945 ;
        RECT 125.090 187.610 128.200 187.805 ;
        RECT 93.370 185.605 94.620 186.655 ;
        RECT 110.640 185.775 111.660 186.835 ;
        RECT 48.720 183.320 50.990 185.270 ;
        RECT 48.800 176.975 52.490 181.625 ;
        RECT 0.950 174.490 8.390 174.950 ;
        RECT 125.090 174.490 128.090 187.610 ;
        RECT 136.280 180.625 137.910 189.480 ;
        RECT 132.600 178.135 138.040 180.625 ;
        RECT 143.720 175.095 144.220 178.465 ;
        RECT 147.400 175.045 148.020 178.605 ;
        RECT 0.950 171.490 128.180 174.490 ;
        RECT 0.950 170.590 8.390 171.490 ;
        RECT 36.545 158.835 83.860 160.445 ;
        RECT 0.960 148.895 11.860 153.515 ;
        RECT 0.960 30.385 5.130 33.865 ;
        RECT 36.545 9.405 38.155 158.835 ;
        RECT 40.740 155.345 42.140 155.350 ;
        RECT 40.540 153.895 47.680 155.345 ;
        RECT 40.740 28.830 42.140 153.895 ;
        RECT 51.730 147.115 55.840 149.355 ;
        RECT 82.250 137.555 83.860 158.835 ;
        RECT 101.810 150.565 103.170 151.925 ;
        RECT 85.220 147.400 86.750 147.410 ;
        RECT 85.050 144.900 87.090 147.400 ;
        RECT 85.100 144.885 87.000 144.900 ;
        RECT 82.200 134.825 83.860 137.555 ;
        RECT 85.220 131.295 87.000 144.885 ;
        RECT 88.260 141.570 88.670 141.945 ;
        RECT 98.350 141.570 99.390 141.585 ;
        RECT 88.260 141.100 99.390 141.570 ;
        RECT 88.260 141.065 88.670 141.100 ;
        RECT 98.350 141.085 99.390 141.100 ;
        RECT 91.200 139.390 92.370 140.595 ;
        RECT 91.200 139.265 99.260 139.390 ;
        RECT 91.200 139.145 99.360 139.265 ;
        RECT 91.270 138.720 99.360 139.145 ;
        RECT 97.790 138.615 99.360 138.720 ;
        RECT 104.990 135.100 128.850 165.500 ;
        RECT 130.050 135.100 153.910 165.500 ;
        RECT 111.450 132.050 115.270 134.660 ;
        RECT 111.530 131.995 114.420 132.050 ;
        RECT 81.360 128.535 83.600 131.115 ;
        RECT 85.170 129.745 87.620 131.295 ;
        RECT 108.720 129.755 111.090 131.345 ;
        RECT 111.530 126.170 114.390 131.995 ;
        RECT 139.990 126.170 145.120 126.200 ;
        RECT 81.300 126.140 145.120 126.170 ;
        RECT 81.040 125.510 145.120 126.140 ;
        RECT 81.040 125.500 144.950 125.510 ;
        RECT 81.040 125.460 85.150 125.500 ;
        RECT 51.240 95.800 81.700 125.000 ;
        RECT 82.900 95.800 113.360 125.000 ;
        RECT 114.560 95.800 145.020 125.000 ;
        RECT 51.240 65.400 81.700 94.600 ;
        RECT 82.900 65.400 113.360 94.600 ;
        RECT 114.560 65.400 145.020 94.600 ;
        RECT 51.240 35.000 81.700 64.200 ;
        RECT 82.900 35.000 113.360 64.200 ;
        RECT 114.560 35.000 145.020 64.200 ;
        RECT 143.690 30.345 144.280 32.765 ;
        RECT 147.300 30.285 148.060 32.745 ;
        RECT 40.740 27.220 69.255 28.830 ;
        RECT 40.740 27.030 42.140 27.220 ;
        RECT 67.645 13.960 69.255 27.220 ;
        RECT 136.790 22.985 138.260 24.505 ;
        RECT 126.820 18.485 128.480 20.265 ;
        RECT 96.580 17.035 98.930 18.175 ;
        RECT 147.210 15.395 148.350 16.605 ;
        RECT 155.780 15.950 157.090 16.465 ;
        RECT 155.250 15.350 159.120 15.950 ;
        RECT 155.780 15.085 157.090 15.350 ;
        RECT 40.780 9.405 47.040 9.500 ;
        RECT 36.545 7.795 47.040 9.405 ;
        RECT 40.780 7.770 47.040 7.795 ;
        RECT 48.920 5.155 52.990 7.435 ;
        RECT 67.570 5.310 69.510 13.960 ;
        RECT 146.930 10.895 148.090 12.305 ;
        RECT 152.785 5.390 153.375 5.415 ;
        RECT 158.520 5.390 159.120 15.350 ;
        RECT 67.645 5.245 69.255 5.310 ;
        RECT 152.780 4.790 159.120 5.390 ;
        RECT 152.785 4.765 153.375 4.790 ;
      LAYER met4 ;
        RECT 3.990 223.990 4.290 224.760 ;
        RECT 7.670 223.990 7.970 224.760 ;
        RECT 3.990 223.690 7.970 223.990 ;
        RECT 3.990 222.915 4.290 223.690 ;
        RECT 3.975 222.585 4.305 222.915 ;
        RECT 11.350 220.470 11.650 224.760 ;
        RECT 15.030 220.470 15.330 224.760 ;
        RECT 16.795 220.470 17.125 220.485 ;
        RECT 2.500 220.170 17.125 220.470 ;
        RECT 16.795 220.155 17.125 220.170 ;
        RECT 18.710 219.120 19.010 224.760 ;
        RECT 22.390 219.145 22.690 224.760 ;
        RECT 26.070 221.225 26.370 224.760 ;
        RECT 26.045 220.095 26.415 221.225 ;
        RECT 29.750 220.130 30.050 224.760 ;
        RECT 40.790 221.250 41.090 224.760 ;
        RECT 44.470 221.670 44.770 224.760 ;
        RECT 55.510 222.510 55.810 224.760 ;
        RECT 60.745 222.510 62.005 222.535 ;
        RECT 55.510 222.210 62.005 222.510 ;
        RECT 60.745 222.205 62.005 222.210 ;
        RECT 44.390 221.370 55.840 221.670 ;
        RECT 40.790 221.075 41.120 221.250 ;
        RECT 40.565 220.705 42.405 221.075 ;
        RECT 49.000 220.760 50.500 220.770 ;
        RECT 29.750 219.830 49.000 220.130 ;
        RECT 54.155 219.875 54.495 220.775 ;
        RECT 55.540 220.265 55.840 221.370 ;
        RECT 62.870 221.215 63.170 224.760 ;
        RECT 66.550 223.165 66.850 224.760 ;
        RECT 70.230 224.625 70.530 224.760 ;
        RECT 68.225 224.440 70.530 224.625 ;
        RECT 68.225 224.115 70.525 224.440 ;
        RECT 73.910 223.870 74.210 224.760 ;
        RECT 71.690 223.410 74.260 223.870 ;
        RECT 77.590 223.450 77.890 224.760 ;
        RECT 81.270 224.280 81.570 224.760 ;
        RECT 83.095 224.280 83.425 224.295 ;
        RECT 81.270 223.980 83.425 224.280 ;
        RECT 83.095 223.965 83.425 223.980 ;
        RECT 79.365 223.450 79.695 223.465 ;
        RECT 65.175 222.835 67.375 223.165 ;
        RECT 77.590 223.150 79.695 223.450 ;
        RECT 79.365 223.135 79.695 223.150 ;
        RECT 64.215 222.490 65.705 222.535 ;
        RECT 64.215 222.190 80.900 222.490 ;
        RECT 64.215 222.185 65.705 222.190 ;
        RECT 60.835 220.885 63.255 221.215 ;
        RECT 62.870 220.830 63.170 220.885 ;
        RECT 22.375 219.120 22.705 219.145 ;
        RECT 18.710 218.820 22.810 219.120 ;
        RECT 22.375 218.815 22.705 218.820 ;
        RECT 48.995 218.115 49.000 219.365 ;
        RECT 50.500 218.115 50.535 219.365 ;
        RECT 48.775 212.045 49.000 214.535 ;
        RECT 50.500 212.045 50.875 214.535 ;
        RECT 54.190 212.895 54.490 219.875 ;
        RECT 55.005 218.635 56.145 220.265 ;
        RECT 54.190 212.060 55.615 212.895 ;
        RECT 54.205 211.835 55.615 212.060 ;
        RECT 78.875 211.350 79.205 211.680 ;
        RECT 9.035 209.120 12.405 209.195 ;
        RECT 42.645 209.120 45.155 209.125 ;
        RECT 2.500 206.620 45.290 209.120 ;
        RECT 9.035 206.435 12.405 206.620 ;
        RECT 42.645 206.615 45.155 206.620 ;
        RECT 43.500 206.610 45.000 206.615 ;
        RECT 48.990 206.565 49.000 209.165 ;
        RECT 50.500 206.565 50.510 209.165 ;
        RECT 75.295 206.675 78.395 209.115 ;
        RECT 50.500 199.555 52.575 202.095 ;
        RECT 78.890 195.360 79.190 211.350 ;
        RECT 79.795 210.615 80.125 210.945 ;
        RECT 79.810 196.725 80.110 210.615 ;
        RECT 80.600 206.240 80.900 222.190 ;
        RECT 84.950 210.905 85.250 224.760 ;
        RECT 88.630 211.760 88.930 224.760 ;
        RECT 88.560 211.320 89.040 211.760 ;
        RECT 92.310 211.265 92.610 224.760 ;
        RECT 95.990 211.875 96.290 224.760 ;
        RECT 107.030 213.505 107.330 224.760 ;
        RECT 110.710 219.465 111.010 224.760 ;
        RECT 109.815 218.915 111.205 219.465 ;
        RECT 106.575 212.365 107.675 213.505 ;
        RECT 95.895 211.285 96.455 211.875 ;
        RECT 84.935 210.575 85.265 210.905 ;
        RECT 92.295 210.345 93.025 211.265 ;
        RECT 80.600 205.940 85.270 206.240 ;
        RECT 84.605 203.725 85.250 205.940 ;
        RECT 118.070 204.705 118.370 224.760 ;
        RECT 119.770 211.925 120.070 211.940 ;
        RECT 119.675 211.335 120.235 211.925 ;
        RECT 119.680 211.320 120.210 211.335 ;
        RECT 84.950 203.590 85.250 203.725 ;
        RECT 117.045 203.625 118.385 204.705 ;
        RECT 118.070 203.590 118.370 203.625 ;
        RECT 79.775 196.265 80.165 196.725 ;
        RECT 94.325 195.360 95.335 195.515 ;
        RECT 78.890 195.060 95.335 195.360 ;
        RECT 94.180 194.870 95.335 195.060 ;
        RECT 94.325 194.505 95.335 194.870 ;
        RECT 110.755 195.050 111.635 195.545 ;
        RECT 119.910 195.050 120.210 211.320 ;
        RECT 120.935 210.305 122.005 210.835 ;
        RECT 110.755 194.750 120.240 195.050 ;
        RECT 110.755 194.415 111.635 194.750 ;
        RECT 79.690 193.610 80.320 194.180 ;
        RECT 79.775 186.405 80.110 193.610 ;
        RECT 93.415 186.405 94.425 186.635 ;
        RECT 79.775 186.045 94.425 186.405 ;
        RECT 79.775 186.040 80.075 186.045 ;
        RECT 93.415 185.625 94.425 186.045 ;
        RECT 110.685 186.460 111.615 186.815 ;
        RECT 121.500 186.460 121.800 210.305 ;
        RECT 125.430 191.740 125.730 224.760 ;
        RECT 132.790 224.410 133.090 224.760 ;
        RECT 128.185 222.385 128.765 223.465 ;
        RECT 129.505 223.325 130.115 224.285 ;
        RECT 131.160 224.110 133.090 224.410 ;
        RECT 128.460 217.065 128.760 222.385 ;
        RECT 128.455 216.295 129.225 217.065 ;
        RECT 128.460 216.250 128.760 216.295 ;
        RECT 129.810 208.540 130.110 223.325 ;
        RECT 131.160 211.385 131.460 224.110 ;
        RECT 136.470 222.075 136.770 224.760 ;
        RECT 136.455 221.745 136.785 222.075 ;
        RECT 140.150 222.015 140.450 224.760 ;
        RECT 140.025 219.215 140.635 222.015 ;
        RECT 130.995 209.645 131.715 211.385 ;
        RECT 131.160 209.620 131.460 209.645 ;
        RECT 129.810 208.225 130.140 208.540 ;
        RECT 129.810 206.185 130.955 208.225 ;
        RECT 129.810 206.140 130.110 206.185 ;
        RECT 123.020 191.440 125.730 191.740 ;
        RECT 110.685 186.160 121.800 186.460 ;
        RECT 110.685 185.795 111.615 186.160 ;
        RECT 48.765 183.315 49.000 185.275 ;
        RECT 50.500 183.315 50.945 185.275 ;
        RECT 50.500 176.995 52.445 181.605 ;
        RECT 0.995 170.585 1.000 174.955 ;
        RECT 2.500 170.585 8.345 174.955 ;
        RECT 123.025 169.665 123.325 191.440 ;
        RECT 143.830 178.445 144.130 224.760 ;
        RECT 147.810 224.750 147.815 225.750 ;
        RECT 147.510 178.585 147.815 224.750 ;
        RECT 143.765 175.115 144.175 178.445 ;
        RECT 147.445 175.065 147.975 178.585 ;
        RECT 54.315 169.365 123.325 169.665 ;
        RECT 2.500 148.915 11.815 153.495 ;
        RECT 54.315 149.335 54.615 169.365 ;
        RECT 101.870 166.070 134.630 167.030 ;
        RECT 101.870 152.860 102.830 166.070 ;
        RECT 114.880 165.105 115.840 166.070 ;
        RECT 101.800 150.580 103.160 152.860 ;
        RECT 101.860 150.510 103.120 150.580 ;
        RECT 51.775 147.135 55.795 149.335 ;
        RECT 101.860 147.480 103.010 150.510 ;
        RECT 85.340 147.405 104.630 147.480 ;
        RECT 85.095 144.970 104.630 147.405 ;
        RECT 85.095 144.895 87.045 144.970 ;
        RECT 105.385 135.495 126.995 165.105 ;
        RECT 128.350 135.200 128.830 165.440 ;
        RECT 133.670 165.105 134.630 166.070 ;
        RECT 130.445 135.495 152.055 165.105 ;
        RECT 153.410 135.380 153.890 165.440 ;
        RECT 111.495 134.550 115.225 134.665 ;
        RECT 111.495 133.965 116.510 134.550 ;
        RECT 128.350 133.965 128.960 135.200 ;
        RECT 153.410 135.160 154.300 135.380 ;
        RECT 153.460 133.965 154.300 135.160 ;
        RECT 111.495 132.760 154.300 133.965 ;
        RECT 111.495 132.675 154.115 132.760 ;
        RECT 111.495 132.045 116.510 132.675 ;
        RECT 115.060 131.870 116.510 132.045 ;
        RECT 108.765 131.280 111.045 131.325 ;
        RECT 81.405 130.490 83.555 131.095 ;
        RECT 50.500 128.600 83.555 130.490 ;
        RECT 108.765 129.775 111.060 131.280 ;
        RECT 81.405 128.555 83.555 128.600 ;
        RECT 108.850 127.800 111.060 129.775 ;
        RECT 65.480 126.550 129.360 127.800 ;
        RECT 65.480 124.605 66.000 126.550 ;
        RECT 81.085 125.455 85.105 126.145 ;
        RECT 51.635 96.195 79.845 124.605 ;
        RECT 65.480 94.205 66.000 96.195 ;
        RECT 51.635 65.795 79.845 94.205 ;
        RECT 65.480 63.805 66.000 65.795 ;
        RECT 51.635 35.395 79.845 63.805 ;
        RECT 65.480 34.400 66.000 35.395 ;
        RECT 81.180 34.400 81.700 125.455 ;
        RECT 97.140 124.605 97.660 126.550 ;
        RECT 110.775 125.495 115.165 126.175 ;
        RECT 83.295 96.195 111.505 124.605 ;
        RECT 97.140 94.205 97.660 96.195 ;
        RECT 83.295 65.795 111.505 94.205 ;
        RECT 97.140 63.805 97.660 65.795 ;
        RECT 83.295 35.395 111.505 63.805 ;
        RECT 97.140 34.400 97.660 35.395 ;
        RECT 112.840 34.400 113.360 125.495 ;
        RECT 128.800 124.605 129.320 126.550 ;
        RECT 140.035 125.505 145.075 126.205 ;
        RECT 114.955 96.195 143.165 124.605 ;
        RECT 128.800 94.205 129.320 96.195 ;
        RECT 114.955 65.795 143.165 94.205 ;
        RECT 128.800 63.805 129.320 65.795 ;
        RECT 114.955 35.395 143.165 63.805 ;
        RECT 128.800 34.400 129.320 35.395 ;
        RECT 144.500 34.400 145.020 125.505 ;
        RECT 2.500 30.405 5.085 33.845 ;
        RECT 143.735 30.365 144.235 32.745 ;
        RECT 147.515 32.725 147.815 32.730 ;
        RECT 136.835 24.040 138.215 24.485 ;
        RECT 134.670 23.440 138.215 24.040 ;
        RECT 126.865 18.505 128.435 20.245 ;
        RECT 96.625 17.650 98.885 18.155 ;
        RECT 90.320 17.055 98.885 17.650 ;
        RECT 90.320 17.050 98.770 17.055 ;
        RECT 40.825 7.765 46.995 9.505 ;
        RECT 46.160 1.000 46.760 7.765 ;
        RECT 50.500 5.175 52.945 7.415 ;
        RECT 67.615 5.305 69.465 13.965 ;
        RECT 68.240 1.000 68.840 5.305 ;
        RECT 90.320 1.000 90.920 17.050 ;
        RECT 127.260 4.440 127.860 18.505 ;
        RECT 134.670 8.960 135.270 23.440 ;
        RECT 136.835 23.005 138.215 23.440 ;
        RECT 143.830 12.090 144.130 30.365 ;
        RECT 147.345 30.305 148.015 32.725 ;
        RECT 147.515 16.585 147.815 30.305 ;
        RECT 147.255 15.415 148.305 16.585 ;
        RECT 146.975 12.090 148.045 12.285 ;
        RECT 143.830 11.790 148.045 12.090 ;
        RECT 146.975 10.915 148.045 11.790 ;
        RECT 156.560 8.960 157.160 9.000 ;
        RECT 134.670 8.360 157.200 8.960 ;
        RECT 134.670 8.300 135.270 8.360 ;
        RECT 112.400 3.840 127.860 4.440 ;
        RECT 134.480 4.790 153.380 5.390 ;
        RECT 112.400 1.000 113.000 3.840 ;
        RECT 134.480 1.000 135.080 4.790 ;
        RECT 156.560 1.000 157.160 8.360 ;
  END
END tt_um_vks_pll
END LIBRARY

