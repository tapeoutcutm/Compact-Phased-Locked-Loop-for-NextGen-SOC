magic
tech sky130A
magscale 1 2
timestamp 1712816020
<< locali >>
rect 6280 -1445 6500 -1426
rect 4552 -1656 4948 -1650
rect 4552 -1762 4553 -1656
rect 4947 -1762 4948 -1656
rect 6280 -1695 6301 -1445
rect 6479 -1468 6500 -1445
rect 6479 -1695 6634 -1468
rect 6280 -1714 6634 -1695
rect 4552 -1768 4948 -1762
rect 4646 -1816 4896 -1768
rect 4272 -1974 4896 -1816
rect 6500 -1898 6634 -1714
rect 4272 -2088 4900 -1974
rect 4648 -2096 4900 -2088
rect 6122 -3896 6332 -3500
rect 4094 -4396 4250 -4364
rect 4094 -4452 4240 -4396
rect 3350 -4536 3474 -4460
rect 4092 -4464 4240 -4452
rect 4288 -4464 4380 -4456
rect 4092 -4470 4380 -4464
rect 4092 -4504 4317 -4470
rect 4351 -4504 4380 -4470
rect 4092 -4518 4380 -4504
rect 3350 -4568 3510 -4536
rect 4092 -4538 4348 -4518
rect 4092 -4540 4210 -4538
rect 3350 -4587 3632 -4568
rect 4766 -4584 4880 -4492
rect 3350 -4604 3516 -4587
rect 3344 -4692 3516 -4604
rect 3506 -4693 3516 -4692
rect 3622 -4693 3632 -4587
rect 3506 -4712 3632 -4693
rect 4704 -4587 4920 -4584
rect 4704 -4693 4723 -4587
rect 4901 -4693 4920 -4587
rect 4704 -4696 4920 -4693
rect 5072 -4709 5698 -4674
rect 5072 -4743 5104 -4709
rect 5138 -4743 5698 -4709
rect 5072 -4778 5698 -4743
rect 5112 -4794 5698 -4778
<< viali >>
rect 4553 -1762 4947 -1656
rect 6301 -1695 6479 -1445
rect 4317 -4504 4351 -4470
rect 3516 -4693 3622 -4587
rect 4723 -4693 4901 -4587
rect 5104 -4743 5138 -4709
<< metal1 >>
rect 4794 -1355 5054 -1354
rect 4794 -1599 4834 -1355
rect 5014 -1599 5054 -1355
rect 4794 -1600 5054 -1599
rect 6274 -1445 6506 -1414
rect 4540 -1656 4960 -1644
rect 4540 -1762 4553 -1656
rect 4947 -1762 4960 -1656
rect 6274 -1695 6301 -1445
rect 6479 -1695 6506 -1445
rect 6274 -1702 6332 -1695
rect 6448 -1702 6506 -1695
rect 6274 -1726 6506 -1702
rect 4540 -1774 4960 -1762
rect 6040 -1870 6422 -1866
rect 3590 -1882 4180 -1876
rect 3520 -1952 4180 -1882
rect 6040 -1904 6532 -1870
rect 3520 -2468 3674 -1952
rect 5294 -1968 5374 -1962
rect 5018 -2028 5374 -1968
rect 3912 -2074 4012 -2068
rect 3912 -2126 3936 -2074
rect 3988 -2126 4012 -2074
rect 3912 -2138 4012 -2126
rect 3912 -2190 3936 -2138
rect 3988 -2190 4012 -2138
rect 3912 -2202 4012 -2190
rect 3912 -2254 3936 -2202
rect 3988 -2254 4012 -2202
rect 3912 -2266 4012 -2254
rect 3912 -2318 3936 -2266
rect 3988 -2318 4012 -2266
rect 3912 -2324 4012 -2318
rect 4144 -2076 4244 -2070
rect 4144 -2128 4168 -2076
rect 4220 -2128 4244 -2076
rect 4144 -2140 4244 -2128
rect 4144 -2192 4168 -2140
rect 4220 -2192 4244 -2140
rect 4144 -2204 4244 -2192
rect 4144 -2256 4168 -2204
rect 4220 -2256 4244 -2204
rect 5064 -2109 5172 -2106
rect 5064 -2161 5092 -2109
rect 5144 -2161 5172 -2109
rect 5064 -2173 5172 -2161
rect 5064 -2225 5092 -2173
rect 5144 -2225 5172 -2173
rect 5064 -2228 5172 -2225
rect 5294 -2108 5374 -2028
rect 6040 -2108 6112 -1904
rect 4144 -2268 4244 -2256
rect 4144 -2320 4168 -2268
rect 4220 -2320 4244 -2268
rect 4144 -2326 4244 -2320
rect 3470 -2476 3674 -2468
rect 3294 -2676 3674 -2476
rect 3470 -2698 3674 -2676
rect 3520 -3234 3674 -2698
rect 5294 -2434 5364 -2108
rect 6042 -2434 6112 -2108
rect 6328 -2068 6416 -2048
rect 6328 -2120 6346 -2068
rect 6398 -2120 6416 -2068
rect 6328 -2132 6416 -2120
rect 6328 -2184 6346 -2132
rect 6398 -2184 6416 -2132
rect 6328 -2196 6416 -2184
rect 6328 -2248 6346 -2196
rect 6398 -2248 6416 -2196
rect 6328 -2268 6416 -2248
rect 3786 -2878 3902 -2852
rect 3786 -2930 3818 -2878
rect 3870 -2930 3902 -2878
rect 3786 -2942 3902 -2930
rect 3786 -2994 3818 -2942
rect 3870 -2994 3902 -2942
rect 3786 -3006 3902 -2994
rect 3786 -3058 3818 -3006
rect 3870 -3058 3902 -3006
rect 3786 -3070 3902 -3058
rect 3786 -3122 3818 -3070
rect 3870 -3122 3902 -3070
rect 3786 -3148 3902 -3122
rect 4030 -2884 4146 -2858
rect 4030 -2936 4062 -2884
rect 4114 -2936 4146 -2884
rect 4030 -2948 4146 -2936
rect 4030 -3000 4062 -2948
rect 4114 -3000 4146 -2948
rect 4030 -3012 4146 -3000
rect 4030 -3064 4062 -3012
rect 4114 -3064 4146 -3012
rect 5294 -3020 6112 -2434
rect 5294 -3046 5376 -3020
rect 4030 -3076 4146 -3064
rect 4030 -3128 4062 -3076
rect 4114 -3128 4146 -3076
rect 4030 -3154 4146 -3128
rect 4790 -3204 5018 -3062
rect 3520 -3284 4150 -3234
rect 3532 -3304 4150 -3284
rect 4222 -3489 4376 -3474
rect 4222 -3605 4241 -3489
rect 4357 -3494 4376 -3489
rect 4790 -3490 4976 -3204
rect 5294 -3298 5370 -3046
rect 5024 -3352 5370 -3298
rect 5024 -3358 5348 -3352
rect 5548 -3372 5856 -3020
rect 6054 -3346 6112 -3020
rect 6216 -3063 6310 -3048
rect 6216 -3115 6237 -3063
rect 6289 -3115 6310 -3063
rect 6216 -3127 6310 -3115
rect 6216 -3179 6237 -3127
rect 6289 -3179 6310 -3127
rect 6216 -3191 6310 -3179
rect 6216 -3243 6237 -3191
rect 6289 -3243 6310 -3191
rect 6216 -3258 6310 -3243
rect 6446 -3067 6540 -3052
rect 6446 -3119 6467 -3067
rect 6519 -3119 6540 -3067
rect 6446 -3131 6540 -3119
rect 6446 -3183 6467 -3131
rect 6519 -3183 6540 -3131
rect 6446 -3195 6540 -3183
rect 6446 -3247 6467 -3195
rect 6519 -3247 6540 -3195
rect 6446 -3262 6540 -3247
rect 6048 -3372 6112 -3346
rect 5548 -3384 5860 -3372
rect 5552 -3490 5860 -3384
rect 6040 -3394 6112 -3372
rect 6040 -3454 6478 -3394
rect 4790 -3494 5860 -3490
rect 4357 -3605 5860 -3494
rect 4222 -3620 5860 -3605
rect 4790 -3626 4976 -3620
rect 3986 -3716 4078 -3710
rect 4152 -3716 4388 -3712
rect 3986 -3718 4388 -3716
rect 4558 -3718 4614 -3716
rect 3590 -3791 3758 -3790
rect 3590 -3808 3616 -3791
rect 3518 -3820 3616 -3808
rect 3508 -3834 3616 -3820
rect 3506 -3843 3616 -3834
rect 3668 -3843 3680 -3791
rect 3732 -3808 3758 -3791
rect 3986 -3796 4614 -3718
rect 3986 -3798 4152 -3796
rect 3986 -3808 4078 -3798
rect 4388 -3800 4614 -3796
rect 3732 -3843 4078 -3808
rect 3506 -3884 4078 -3843
rect 3668 -3892 4078 -3884
rect 3432 -3975 3530 -3944
rect 3432 -4027 3455 -3975
rect 3507 -4027 3530 -3975
rect 3432 -4058 3530 -4027
rect 3538 -4203 3664 -4180
rect 3538 -4255 3575 -4203
rect 3627 -4255 3664 -4203
rect 3538 -4278 3664 -4255
rect 3800 -4256 4078 -3892
rect 4156 -3864 4298 -3848
rect 4156 -3980 4169 -3864
rect 4285 -3980 4298 -3864
rect 4156 -3996 4298 -3980
rect 4558 -3880 4614 -3800
rect 4290 -4105 4438 -4076
rect 4290 -4157 4306 -4105
rect 4358 -4157 4370 -4105
rect 4422 -4157 4438 -4105
rect 4290 -4186 4438 -4157
rect 4558 -4114 4698 -3880
rect 5632 -3906 5818 -3902
rect 5632 -3990 6276 -3906
rect 5646 -3992 6276 -3990
rect 5646 -4044 5828 -3992
rect 4558 -4182 5012 -4114
rect 5356 -4180 5828 -4044
rect 6072 -4154 6176 -4140
rect 3800 -4264 4324 -4256
rect 4558 -4264 4698 -4182
rect 3800 -4338 4698 -4264
rect 4836 -4257 4938 -4236
rect 5356 -4244 5856 -4180
rect 6072 -4206 6098 -4154
rect 6150 -4206 6176 -4154
rect 6072 -4220 6176 -4206
rect 6516 -4218 6537 -4038
rect 6653 -4218 6674 -4038
rect 6834 -4196 7098 -4052
rect 4836 -4309 4861 -4257
rect 4913 -4309 4938 -4257
rect 4836 -4330 4938 -4309
rect 5022 -4279 5160 -4258
rect 5586 -4262 5856 -4244
rect 3800 -4340 4078 -4338
rect 3798 -4344 4078 -4340
rect 3798 -4352 4020 -4344
rect 4312 -4346 4698 -4338
rect 3798 -4354 3826 -4352
rect 4606 -4354 4698 -4346
rect 5022 -4331 5033 -4279
rect 5085 -4331 5097 -4279
rect 5149 -4331 5160 -4279
rect 5022 -4352 5160 -4331
rect 5632 -4276 5856 -4262
rect 6806 -4222 7098 -4196
rect 6806 -4274 6833 -4222
rect 6885 -4274 6897 -4222
rect 6949 -4274 6961 -4222
rect 7013 -4274 7098 -4222
rect 5632 -4308 6284 -4276
rect 6806 -4298 7098 -4274
rect 6806 -4300 7040 -4298
rect 5632 -4332 6314 -4308
rect 3506 -4400 3826 -4354
rect 3520 -4416 3826 -4400
rect 4650 -4394 4698 -4354
rect 5648 -4356 6314 -4332
rect 5656 -4360 6314 -4356
rect 4650 -4410 4990 -4394
rect 6284 -4398 6314 -4360
rect 4276 -4464 4392 -4450
rect 4650 -4462 5016 -4410
rect 4276 -4516 4312 -4464
rect 4364 -4516 4392 -4464
rect 4276 -4524 4392 -4516
rect 5256 -4503 5428 -4500
rect 4300 -4526 4376 -4524
rect 4420 -4554 4524 -4546
rect 3500 -4584 3638 -4556
rect 3500 -4587 3551 -4584
rect 3603 -4587 3638 -4584
rect 3500 -4693 3516 -4587
rect 3622 -4693 3638 -4587
rect 4150 -4566 4240 -4562
rect 4420 -4566 4439 -4554
rect 4150 -4606 4439 -4566
rect 4491 -4606 4524 -4554
rect 4150 -4616 4524 -4606
rect 4692 -4587 4932 -4578
rect 4150 -4618 4462 -4616
rect 4150 -4634 4247 -4618
rect 3500 -4700 3551 -4693
rect 3603 -4700 3638 -4693
rect 3500 -4724 3638 -4700
rect 4192 -4734 4247 -4634
rect 4427 -4722 4462 -4618
rect 4692 -4693 4723 -4587
rect 4901 -4693 4932 -4587
rect 5256 -4619 5284 -4503
rect 5400 -4530 5428 -4503
rect 6842 -4530 6974 -4510
rect 5400 -4619 6974 -4530
rect 5256 -4622 6974 -4619
rect 4692 -4702 4932 -4693
rect 5066 -4703 5176 -4662
rect 4427 -4734 4524 -4722
rect 4192 -4744 4524 -4734
rect 4158 -4746 4524 -4744
rect 4158 -4798 4183 -4746
rect 4235 -4794 4439 -4746
rect 4235 -4798 4246 -4794
rect 4158 -4802 4246 -4798
rect 4426 -4798 4439 -4794
rect 4491 -4798 4524 -4746
rect 5066 -4755 5094 -4703
rect 5146 -4755 5176 -4703
rect 5066 -4790 5176 -4755
rect 5378 -4776 5980 -4708
rect 4426 -4806 4524 -4798
rect 5360 -4796 5980 -4776
rect 5360 -4826 5590 -4796
rect 5360 -4830 5564 -4826
rect 5364 -4998 5564 -4830
rect 5734 -4896 5854 -4878
rect 5734 -4948 5768 -4896
rect 5820 -4948 5854 -4896
rect 5734 -4966 5854 -4948
rect 5362 -5064 5576 -4998
rect 6842 -5008 6974 -4622
rect 5362 -5078 5986 -5064
rect 5384 -5152 5986 -5078
<< via1 >>
rect 4834 -1599 5014 -1355
rect 4612 -1729 4664 -1677
rect 4676 -1729 4728 -1677
rect 4740 -1729 4792 -1677
rect 4804 -1729 4856 -1677
rect 4868 -1729 4920 -1677
rect 6332 -1695 6448 -1458
rect 6332 -1702 6448 -1695
rect 3936 -2126 3988 -2074
rect 3936 -2190 3988 -2138
rect 3936 -2254 3988 -2202
rect 3936 -2318 3988 -2266
rect 4168 -2128 4220 -2076
rect 4168 -2192 4220 -2140
rect 4168 -2256 4220 -2204
rect 5092 -2161 5144 -2109
rect 5092 -2225 5144 -2173
rect 4168 -2320 4220 -2268
rect 6346 -2120 6398 -2068
rect 6346 -2184 6398 -2132
rect 6346 -2248 6398 -2196
rect 3818 -2930 3870 -2878
rect 3818 -2994 3870 -2942
rect 3818 -3058 3870 -3006
rect 3818 -3122 3870 -3070
rect 4062 -2936 4114 -2884
rect 4062 -3000 4114 -2948
rect 4062 -3064 4114 -3012
rect 4062 -3128 4114 -3076
rect 4241 -3605 4357 -3489
rect 6237 -3115 6289 -3063
rect 6237 -3179 6289 -3127
rect 6237 -3243 6289 -3191
rect 6467 -3119 6519 -3067
rect 6467 -3183 6519 -3131
rect 6467 -3247 6519 -3195
rect 3616 -3843 3668 -3791
rect 3680 -3843 3732 -3791
rect 3455 -4027 3507 -3975
rect 3575 -4255 3627 -4203
rect 4169 -3980 4285 -3864
rect 4306 -4157 4358 -4105
rect 4370 -4157 4422 -4105
rect 6098 -4206 6150 -4154
rect 6537 -4218 6653 -4038
rect 4861 -4309 4913 -4257
rect 5033 -4331 5085 -4279
rect 5097 -4331 5149 -4279
rect 6833 -4274 6885 -4222
rect 6897 -4274 6949 -4222
rect 6961 -4274 7013 -4222
rect 4312 -4470 4364 -4464
rect 4312 -4504 4317 -4470
rect 4317 -4504 4351 -4470
rect 4351 -4504 4364 -4470
rect 4312 -4516 4364 -4504
rect 3551 -4587 3603 -4584
rect 3551 -4636 3603 -4587
rect 3551 -4693 3603 -4648
rect 4439 -4606 4491 -4554
rect 3551 -4700 3603 -4693
rect 4247 -4734 4427 -4618
rect 4763 -4660 4815 -4608
rect 4827 -4660 4879 -4608
rect 5284 -4619 5400 -4503
rect 4183 -4798 4235 -4746
rect 4439 -4798 4491 -4746
rect 5094 -4709 5146 -4703
rect 5094 -4743 5104 -4709
rect 5104 -4743 5138 -4709
rect 5138 -4743 5146 -4709
rect 5094 -4755 5146 -4743
rect 5768 -4948 5820 -4896
<< metal2 >>
rect 4732 -1355 5076 -1340
rect 4016 -1472 4258 -1462
rect 4732 -1472 4834 -1355
rect 4016 -1599 4834 -1472
rect 5014 -1472 5076 -1355
rect 6310 -1458 6470 -1440
rect 6310 -1466 6332 -1458
rect 5416 -1472 6332 -1466
rect 5014 -1599 6332 -1472
rect 4016 -1677 6332 -1599
rect 4016 -1724 4612 -1677
rect 4016 -2018 4258 -1724
rect 4600 -1729 4612 -1724
rect 4664 -1729 4676 -1677
rect 4728 -1729 4740 -1677
rect 4792 -1729 4804 -1677
rect 4856 -1729 4868 -1677
rect 4920 -1702 6332 -1677
rect 6448 -1702 6470 -1458
rect 4920 -1720 6470 -1702
rect 4920 -1724 6460 -1720
rect 4920 -1729 4932 -1724
rect 4600 -1758 4932 -1729
rect 3984 -2058 4258 -2018
rect 3922 -2074 4258 -2058
rect 3922 -2078 3936 -2074
rect 3888 -2126 3936 -2078
rect 3988 -2076 4258 -2074
rect 3988 -2126 4168 -2076
rect 3888 -2128 4168 -2126
rect 4220 -2128 4258 -2076
rect 5084 -2096 5258 -1724
rect 5416 -1726 6460 -1724
rect 6256 -1870 6460 -1726
rect 6256 -1872 6462 -1870
rect 3888 -2138 4258 -2128
rect 3888 -2190 3936 -2138
rect 3988 -2140 4258 -2138
rect 3988 -2190 4168 -2140
rect 3888 -2192 4168 -2190
rect 4220 -2192 4258 -2140
rect 3888 -2202 4258 -2192
rect 3888 -2254 3936 -2202
rect 3988 -2204 4258 -2202
rect 3988 -2254 4168 -2204
rect 3888 -2256 4168 -2254
rect 4220 -2256 4258 -2204
rect 5074 -2109 5258 -2096
rect 5074 -2161 5092 -2109
rect 5144 -2161 5258 -2109
rect 5074 -2173 5258 -2161
rect 5074 -2225 5092 -2173
rect 5144 -2198 5258 -2173
rect 6262 -2046 6462 -1872
rect 6262 -2068 6470 -2046
rect 6262 -2120 6346 -2068
rect 6398 -2120 6470 -2068
rect 6262 -2132 6470 -2120
rect 6262 -2184 6346 -2132
rect 6398 -2184 6470 -2132
rect 6262 -2196 6470 -2184
rect 5144 -2225 5162 -2198
rect 5074 -2238 5162 -2225
rect 3888 -2266 4258 -2256
rect 3888 -2316 3936 -2266
rect 3922 -2318 3936 -2316
rect 3988 -2268 4258 -2266
rect 6262 -2248 6346 -2196
rect 6398 -2248 6470 -2196
rect 6262 -2268 6470 -2248
rect 3988 -2318 4168 -2268
rect 3922 -2320 4168 -2318
rect 4220 -2320 4258 -2268
rect 6338 -2278 6406 -2268
rect 3922 -2328 4258 -2320
rect 3922 -2334 4040 -2328
rect 3988 -2338 4040 -2334
rect 4154 -2336 4234 -2328
rect 3796 -2864 3892 -2842
rect 4040 -2864 4136 -2848
rect 3796 -2878 4150 -2864
rect 3796 -2930 3818 -2878
rect 3870 -2884 4150 -2878
rect 3870 -2930 4062 -2884
rect 3796 -2936 4062 -2930
rect 4114 -2936 4150 -2884
rect 3796 -2942 4150 -2936
rect 3796 -2994 3818 -2942
rect 3870 -2948 4150 -2942
rect 3870 -2994 4062 -2948
rect 3796 -3000 4062 -2994
rect 4114 -3000 4150 -2948
rect 3796 -3006 4150 -3000
rect 3796 -3058 3818 -3006
rect 3870 -3012 4150 -3006
rect 3870 -3058 4062 -3012
rect 3796 -3064 4062 -3058
rect 4114 -3064 4150 -3012
rect 3796 -3070 4150 -3064
rect 3796 -3122 3818 -3070
rect 3870 -3076 4150 -3070
rect 3870 -3122 4062 -3076
rect 3796 -3128 4062 -3122
rect 4114 -3128 4150 -3076
rect 3796 -3130 4150 -3128
rect 3716 -3144 4150 -3130
rect 6226 -3063 6300 -3038
rect 6226 -3115 6237 -3063
rect 6289 -3068 6300 -3063
rect 6456 -3067 6530 -3042
rect 6456 -3068 6467 -3067
rect 6289 -3115 6467 -3068
rect 6226 -3119 6467 -3115
rect 6519 -3068 6530 -3067
rect 6519 -3119 6554 -3068
rect 6226 -3127 6554 -3119
rect 3716 -3576 3914 -3144
rect 4040 -3164 4136 -3144
rect 6226 -3179 6237 -3127
rect 6289 -3131 6554 -3127
rect 6289 -3179 6467 -3131
rect 6226 -3183 6467 -3179
rect 6519 -3183 6554 -3131
rect 6226 -3184 6554 -3183
rect 6226 -3191 6642 -3184
rect 6226 -3243 6237 -3191
rect 6289 -3195 6642 -3191
rect 6289 -3243 6467 -3195
rect 6226 -3247 6467 -3243
rect 6519 -3247 6642 -3195
rect 6226 -3254 6642 -3247
rect 6226 -3268 6300 -3254
rect 3294 -3620 3914 -3576
rect 3292 -3680 3914 -3620
rect 4078 -3464 4328 -3460
rect 4078 -3489 4366 -3464
rect 4078 -3605 4241 -3489
rect 4357 -3605 4366 -3489
rect 6406 -3566 6642 -3254
rect 4078 -3630 4366 -3605
rect 3292 -3684 3726 -3680
rect 3292 -3812 3484 -3684
rect 3518 -3690 3726 -3684
rect 3610 -3780 3726 -3690
rect 4078 -3700 4332 -3630
rect 4078 -3706 4258 -3700
rect 3600 -3791 3748 -3780
rect 3292 -3890 3480 -3812
rect 3600 -3843 3616 -3791
rect 3668 -3843 3680 -3791
rect 3732 -3843 3748 -3791
rect 3600 -3854 3748 -3843
rect 4078 -3804 4256 -3706
rect 6410 -3738 6640 -3566
rect 4078 -3838 4258 -3804
rect 4078 -3864 4288 -3838
rect 3292 -3916 3488 -3890
rect 3292 -3934 3516 -3916
rect 3292 -3975 3520 -3934
rect 3292 -4027 3455 -3975
rect 3507 -4027 3520 -3975
rect 4078 -3980 4169 -3864
rect 4285 -3980 4288 -3864
rect 6410 -3920 6644 -3738
rect 4078 -3998 4288 -3980
rect 4866 -3996 4964 -3994
rect 5178 -3996 5312 -3990
rect 4166 -4006 4288 -3998
rect 3292 -4040 3520 -4027
rect 3388 -4048 3520 -4040
rect 3442 -4068 3520 -4048
rect 4300 -4105 4428 -4066
rect 4862 -4082 5312 -3996
rect 4300 -4157 4306 -4105
rect 4358 -4157 4370 -4105
rect 4422 -4118 4428 -4105
rect 4422 -4157 4474 -4118
rect 3544 -4196 3654 -4170
rect 4300 -4196 4474 -4157
rect 3544 -4203 3720 -4196
rect 3544 -4255 3575 -4203
rect 3627 -4254 3720 -4203
rect 3627 -4255 3716 -4254
rect 3544 -4288 3716 -4255
rect 3574 -4574 3716 -4288
rect 4328 -4444 4474 -4196
rect 4866 -4226 4964 -4082
rect 4846 -4246 4964 -4226
rect 4846 -4257 4968 -4246
rect 4846 -4309 4861 -4257
rect 4913 -4309 4968 -4257
rect 4846 -4310 4968 -4309
rect 5032 -4279 5150 -4248
rect 4846 -4340 4928 -4310
rect 5032 -4331 5033 -4279
rect 5085 -4331 5097 -4279
rect 5149 -4331 5150 -4279
rect 5032 -4362 5150 -4331
rect 5032 -4410 5136 -4362
rect 4310 -4446 4474 -4444
rect 4310 -4464 4494 -4446
rect 4310 -4516 4312 -4464
rect 4364 -4516 4494 -4464
rect 4310 -4536 4494 -4516
rect 3542 -4584 3716 -4574
rect 4160 -4566 4230 -4552
rect 4328 -4554 4514 -4536
rect 4328 -4566 4439 -4554
rect 4160 -4584 4439 -4566
rect 3542 -4636 3551 -4584
rect 3603 -4606 4439 -4584
rect 4491 -4578 4514 -4554
rect 4491 -4580 4644 -4578
rect 4491 -4606 4656 -4580
rect 3603 -4618 4656 -4606
rect 3603 -4636 4247 -4618
rect 3542 -4648 4247 -4636
rect 3542 -4700 3551 -4648
rect 3603 -4700 4247 -4648
rect 3542 -4710 4247 -4700
rect 3556 -4734 4247 -4710
rect 4427 -4628 4656 -4618
rect 4746 -4608 4896 -4588
rect 4746 -4628 4763 -4608
rect 4427 -4660 4763 -4628
rect 4815 -4660 4827 -4608
rect 4879 -4628 4896 -4608
rect 5026 -4628 5140 -4410
rect 5178 -4490 5312 -4082
rect 6404 -4028 6640 -3920
rect 6404 -4038 6664 -4028
rect 6082 -4154 6166 -4130
rect 6082 -4206 6098 -4154
rect 6150 -4156 6166 -4154
rect 6150 -4206 6218 -4156
rect 6404 -4202 6537 -4038
rect 6082 -4230 6218 -4206
rect 6526 -4218 6537 -4202
rect 6653 -4218 6664 -4038
rect 6816 -4210 7030 -4186
rect 6526 -4228 6664 -4218
rect 6810 -4222 7030 -4210
rect 6102 -4392 6218 -4230
rect 6810 -4274 6833 -4222
rect 6885 -4274 6897 -4222
rect 6949 -4274 6961 -4222
rect 7013 -4274 7030 -4222
rect 6810 -4310 7030 -4274
rect 6102 -4420 6232 -4392
rect 6810 -4420 6996 -4310
rect 5178 -4503 5418 -4490
rect 5178 -4616 5284 -4503
rect 5266 -4619 5284 -4616
rect 5400 -4619 5418 -4503
rect 5750 -4540 6998 -4420
rect 4879 -4660 5134 -4628
rect 5266 -4632 5418 -4619
rect 5758 -4624 6998 -4540
rect 4427 -4672 5134 -4660
rect 4427 -4703 5148 -4672
rect 4427 -4734 5094 -4703
rect 3556 -4736 5094 -4734
rect 4160 -4746 5094 -4736
rect 4160 -4798 4183 -4746
rect 4235 -4794 4439 -4746
rect 4235 -4798 4236 -4794
rect 4160 -4800 4236 -4798
rect 4168 -4812 4236 -4800
rect 4436 -4798 4439 -4794
rect 4491 -4755 5094 -4746
rect 5146 -4755 5148 -4703
rect 4491 -4756 5148 -4755
rect 4491 -4798 4514 -4756
rect 4626 -4762 4698 -4756
rect 5092 -4786 5148 -4756
rect 4436 -4816 4514 -4798
rect 5760 -4868 5918 -4624
rect 5744 -4896 5918 -4868
rect 5744 -4948 5768 -4896
rect 5820 -4948 5918 -4896
rect 5744 -4954 5918 -4948
rect 5744 -4976 5844 -4954
use sky130_fd_pr__nfet_01v8_PFL2KG  sky130_fd_pr__nfet_01v8_PFL2KG_0
timestamp 1712816020
transform 1 0 4295 0 1 -4027
box -216 -400 216 400
use sky130_fd_pr__pfet_01v8_6QF7WZ  sky130_fd_pr__pfet_01v8_6QF7WZ_0
timestamp 1712816020
transform 1 0 4020 0 1 -2597
box -344 -819 344 819
use sky130_fd_pr__pfet_01v8_VLWSF2  sky130_fd_pr__pfet_01v8_VLWSF2_0
timestamp 1712816020
transform -1 0 6359 0 -1 -4145
box -396 -319 396 319
use sky130_fd_pr__pfet_01v8_6QP7WZ  XM1
timestamp 1712816020
transform 1 0 5052 0 1 -2661
box -226 -819 226 819
use sky130_fd_pr__pfet_01v8_6QN7WZ  XM2
timestamp 1712816020
transform 1 0 6367 0 1 -2651
box -285 -919 285 919
use sky130_fd_pr__nfet_01v8_U4BYG2  XM4
timestamp 1712816020
transform 1 0 6318 0 1 -4932
box -686 -300 686 300
use sky130_fd_pr__nfet_01v8_8PEQNF  XM5
timestamp 1712816020
transform 1 0 4972 0 1 -4290
box -236 -270 236 270
use sky130_fd_pr__nfet_01v8_PFL2KG  XM7
timestamp 1712816020
transform 1 0 3545 0 1 -4119
box -216 -400 216 400
<< labels >>
flabel metal1 s 5364 -5020 5564 -4820 0 FreeSans 626 0 0 0 Qb
port 1 nsew
flabel metal1 s 5356 -4244 5556 -4044 0 FreeSans 626 0 0 0 Qa
port 2 nsew
flabel metal1 s 6884 -4256 7084 -4056 0 FreeSans 626 0 0 0 Vout
port 3 nsew
flabel metal1 s 3294 -2676 3494 -2476 0 FreeSans 626 0 0 0 CP_bias
port 4 nsew
flabel metal2 s 4824 -1580 5024 -1380 0 FreeSans 626 0 0 0 VDD
port 5 nsew
flabel metal2 s 4226 -4784 4426 -4584 0 FreeSans 626 0 0 0 Vss
port 6 nsew
<< end >>
