magic
tech sky130A
magscale 1 2
timestamp 1712816020
<< pwell >>
rect -236 -270 236 270
<< nmos >>
rect -50 -70 50 70
<< ndiff >>
rect -108 51 -50 70
rect -108 17 -96 51
rect -62 17 -50 51
rect -108 -17 -50 17
rect -108 -51 -96 -17
rect -62 -51 -50 -17
rect -108 -70 -50 -51
rect 50 51 108 70
rect 50 17 62 51
rect 96 17 108 51
rect 50 -17 108 17
rect 50 -51 62 -17
rect 96 -51 108 -17
rect 50 -70 108 -51
<< ndiffc >>
rect -96 17 -62 51
rect -96 -51 -62 -17
rect 62 17 96 51
rect 62 -51 96 -17
<< psubdiff >>
rect -210 210 -85 244
rect -51 210 -17 244
rect 17 210 51 244
rect 85 210 210 244
rect -210 119 -176 210
rect -210 51 -176 85
rect 176 119 210 210
rect -210 -17 -176 17
rect -210 -85 -176 -51
rect 176 51 210 85
rect 176 -17 210 17
rect -210 -210 -176 -119
rect 176 -85 210 -51
rect 176 -210 210 -119
rect -210 -244 -85 -210
rect -51 -244 -17 -210
rect 17 -244 51 -210
rect 85 -244 210 -210
<< psubdiffcont >>
rect -85 210 -51 244
rect -17 210 17 244
rect 51 210 85 244
rect -210 85 -176 119
rect 176 85 210 119
rect -210 17 -176 51
rect -210 -51 -176 -17
rect 176 17 210 51
rect 176 -51 210 -17
rect -210 -119 -176 -85
rect 176 -119 210 -85
rect -85 -244 -51 -210
rect -17 -244 17 -210
rect 51 -244 85 -210
<< poly >>
rect -50 142 50 158
rect -50 108 -17 142
rect 17 108 50 142
rect -50 70 50 108
rect -50 -108 50 -70
rect -50 -142 -17 -108
rect 17 -142 50 -108
rect -50 -158 50 -142
<< polycont >>
rect -17 108 17 142
rect -17 -142 17 -108
<< locali >>
rect -210 210 -85 244
rect -51 210 -17 244
rect 17 210 51 244
rect 85 210 210 244
rect -210 119 -176 210
rect -50 108 -17 142
rect 17 108 50 142
rect 176 119 210 210
rect -210 51 -176 85
rect -210 -17 -176 17
rect -210 -85 -176 -51
rect -96 53 -62 74
rect -96 -17 -62 17
rect -96 -74 -62 -53
rect 62 53 96 74
rect 62 -17 96 17
rect 62 -74 96 -53
rect 176 51 210 85
rect 176 -17 210 17
rect 176 -85 210 -51
rect -210 -210 -176 -119
rect -50 -142 -17 -108
rect 17 -142 50 -108
rect 176 -210 210 -119
rect -210 -244 -85 -210
rect -51 -244 -17 -210
rect 17 -244 51 -210
rect 85 -244 210 -210
<< viali >>
rect -17 108 17 142
rect -96 51 -62 53
rect -96 19 -62 51
rect -96 -51 -62 -19
rect -96 -53 -62 -51
rect 62 51 96 53
rect 62 19 96 51
rect 62 -51 96 -19
rect 62 -53 96 -51
rect -17 -142 17 -108
<< metal1 >>
rect -46 142 46 148
rect -46 108 -17 142
rect 17 108 46 142
rect -46 102 46 108
rect -102 53 -56 70
rect -102 19 -96 53
rect -62 19 -56 53
rect -102 -19 -56 19
rect -102 -53 -96 -19
rect -62 -53 -56 -19
rect -102 -70 -56 -53
rect 56 53 102 70
rect 56 19 62 53
rect 96 19 102 53
rect 56 -19 102 19
rect 56 -53 62 -19
rect 96 -53 102 -19
rect 56 -70 102 -53
rect -46 -108 46 -102
rect -46 -142 -17 -108
rect 17 -142 46 -108
rect -46 -148 46 -142
<< properties >>
string FIXED_BBOX -192 -226 192 226
<< end >>
