magic
tech sky130A
magscale 1 2
timestamp 1712816020
<< pwell >>
rect -365 -425 365 425
<< nmos >>
rect -179 -225 -29 225
rect 29 -225 179 225
<< ndiff >>
rect -237 187 -179 225
rect -237 153 -225 187
rect -191 153 -179 187
rect -237 119 -179 153
rect -237 85 -225 119
rect -191 85 -179 119
rect -237 51 -179 85
rect -237 17 -225 51
rect -191 17 -179 51
rect -237 -17 -179 17
rect -237 -51 -225 -17
rect -191 -51 -179 -17
rect -237 -85 -179 -51
rect -237 -119 -225 -85
rect -191 -119 -179 -85
rect -237 -153 -179 -119
rect -237 -187 -225 -153
rect -191 -187 -179 -153
rect -237 -225 -179 -187
rect -29 187 29 225
rect -29 153 -17 187
rect 17 153 29 187
rect -29 119 29 153
rect -29 85 -17 119
rect 17 85 29 119
rect -29 51 29 85
rect -29 17 -17 51
rect 17 17 29 51
rect -29 -17 29 17
rect -29 -51 -17 -17
rect 17 -51 29 -17
rect -29 -85 29 -51
rect -29 -119 -17 -85
rect 17 -119 29 -85
rect -29 -153 29 -119
rect -29 -187 -17 -153
rect 17 -187 29 -153
rect -29 -225 29 -187
rect 179 187 237 225
rect 179 153 191 187
rect 225 153 237 187
rect 179 119 237 153
rect 179 85 191 119
rect 225 85 237 119
rect 179 51 237 85
rect 179 17 191 51
rect 225 17 237 51
rect 179 -17 237 17
rect 179 -51 191 -17
rect 225 -51 237 -17
rect 179 -85 237 -51
rect 179 -119 191 -85
rect 225 -119 237 -85
rect 179 -153 237 -119
rect 179 -187 191 -153
rect 225 -187 237 -153
rect 179 -225 237 -187
<< ndiffc >>
rect -225 153 -191 187
rect -225 85 -191 119
rect -225 17 -191 51
rect -225 -51 -191 -17
rect -225 -119 -191 -85
rect -225 -187 -191 -153
rect -17 153 17 187
rect -17 85 17 119
rect -17 17 17 51
rect -17 -51 17 -17
rect -17 -119 17 -85
rect -17 -187 17 -153
rect 191 153 225 187
rect 191 85 225 119
rect 191 17 225 51
rect 191 -51 225 -17
rect 191 -119 225 -85
rect 191 -187 225 -153
<< psubdiff >>
rect -339 365 -221 399
rect -187 365 -153 399
rect -119 365 -85 399
rect -51 365 -17 399
rect 17 365 51 399
rect 85 365 119 399
rect 153 365 187 399
rect 221 365 339 399
rect -339 289 -305 365
rect -339 221 -305 255
rect 305 289 339 365
rect -339 153 -305 187
rect -339 85 -305 119
rect -339 17 -305 51
rect -339 -51 -305 -17
rect -339 -119 -305 -85
rect -339 -187 -305 -153
rect -339 -255 -305 -221
rect 305 221 339 255
rect 305 153 339 187
rect 305 85 339 119
rect 305 17 339 51
rect 305 -51 339 -17
rect 305 -119 339 -85
rect 305 -187 339 -153
rect -339 -365 -305 -289
rect 305 -255 339 -221
rect 305 -365 339 -289
rect -339 -399 -221 -365
rect -187 -399 -153 -365
rect -119 -399 -85 -365
rect -51 -399 -17 -365
rect 17 -399 51 -365
rect 85 -399 119 -365
rect 153 -399 187 -365
rect 221 -399 339 -365
<< psubdiffcont >>
rect -221 365 -187 399
rect -153 365 -119 399
rect -85 365 -51 399
rect -17 365 17 399
rect 51 365 85 399
rect 119 365 153 399
rect 187 365 221 399
rect -339 255 -305 289
rect 305 255 339 289
rect -339 187 -305 221
rect -339 119 -305 153
rect -339 51 -305 85
rect -339 -17 -305 17
rect -339 -85 -305 -51
rect -339 -153 -305 -119
rect -339 -221 -305 -187
rect 305 187 339 221
rect 305 119 339 153
rect 305 51 339 85
rect 305 -17 339 17
rect 305 -85 339 -51
rect 305 -153 339 -119
rect 305 -221 339 -187
rect -339 -289 -305 -255
rect 305 -289 339 -255
rect -221 -399 -187 -365
rect -153 -399 -119 -365
rect -85 -399 -51 -365
rect -17 -399 17 -365
rect 51 -399 85 -365
rect 119 -399 153 -365
rect 187 -399 221 -365
<< poly >>
rect -179 297 -29 313
rect -179 263 -155 297
rect -121 263 -87 297
rect -53 263 -29 297
rect -179 225 -29 263
rect 29 297 179 313
rect 29 263 53 297
rect 87 263 121 297
rect 155 263 179 297
rect 29 225 179 263
rect -179 -263 -29 -225
rect -179 -297 -155 -263
rect -121 -297 -87 -263
rect -53 -297 -29 -263
rect -179 -313 -29 -297
rect 29 -263 179 -225
rect 29 -297 53 -263
rect 87 -297 121 -263
rect 155 -297 179 -263
rect 29 -313 179 -297
<< polycont >>
rect -155 263 -121 297
rect -87 263 -53 297
rect 53 263 87 297
rect 121 263 155 297
rect -155 -297 -121 -263
rect -87 -297 -53 -263
rect 53 -297 87 -263
rect 121 -297 155 -263
<< locali >>
rect -339 365 -221 399
rect -187 365 -153 399
rect -119 365 -85 399
rect -51 365 -17 399
rect 17 365 51 399
rect 85 365 119 399
rect 153 365 187 399
rect 221 365 339 399
rect -339 289 -305 365
rect -179 263 -157 297
rect -121 263 -87 297
rect -51 263 -29 297
rect 29 263 51 297
rect 87 263 121 297
rect 157 263 179 297
rect 305 289 339 365
rect -339 221 -305 255
rect -339 153 -305 187
rect -339 85 -305 119
rect -339 17 -305 51
rect -339 -51 -305 -17
rect -339 -119 -305 -85
rect -339 -187 -305 -153
rect -339 -255 -305 -221
rect -225 197 -191 229
rect -225 125 -191 153
rect -225 53 -191 85
rect -225 -17 -191 17
rect -225 -85 -191 -53
rect -225 -153 -191 -125
rect -225 -229 -191 -197
rect -17 197 17 229
rect -17 125 17 153
rect -17 53 17 85
rect -17 -17 17 17
rect -17 -85 17 -53
rect -17 -153 17 -125
rect -17 -229 17 -197
rect 191 197 225 229
rect 191 125 225 153
rect 191 53 225 85
rect 191 -17 225 17
rect 191 -85 225 -53
rect 191 -153 225 -125
rect 191 -229 225 -197
rect 305 221 339 255
rect 305 153 339 187
rect 305 85 339 119
rect 305 17 339 51
rect 305 -51 339 -17
rect 305 -119 339 -85
rect 305 -187 339 -153
rect 305 -255 339 -221
rect -339 -365 -305 -289
rect -179 -297 -157 -263
rect -121 -297 -87 -263
rect -51 -297 -29 -263
rect 29 -297 51 -263
rect 87 -297 121 -263
rect 157 -297 179 -263
rect 305 -365 339 -289
rect -339 -399 -221 -365
rect -187 -399 -153 -365
rect -119 -399 -85 -365
rect -51 -399 -17 -365
rect 17 -399 51 -365
rect 85 -399 119 -365
rect 153 -399 187 -365
rect 221 -399 339 -365
<< viali >>
rect -157 263 -155 297
rect -155 263 -123 297
rect -85 263 -53 297
rect -53 263 -51 297
rect 51 263 53 297
rect 53 263 85 297
rect 123 263 155 297
rect 155 263 157 297
rect -225 187 -191 197
rect -225 163 -191 187
rect -225 119 -191 125
rect -225 91 -191 119
rect -225 51 -191 53
rect -225 19 -191 51
rect -225 -51 -191 -19
rect -225 -53 -191 -51
rect -225 -119 -191 -91
rect -225 -125 -191 -119
rect -225 -187 -191 -163
rect -225 -197 -191 -187
rect -17 187 17 197
rect -17 163 17 187
rect -17 119 17 125
rect -17 91 17 119
rect -17 51 17 53
rect -17 19 17 51
rect -17 -51 17 -19
rect -17 -53 17 -51
rect -17 -119 17 -91
rect -17 -125 17 -119
rect -17 -187 17 -163
rect -17 -197 17 -187
rect 191 187 225 197
rect 191 163 225 187
rect 191 119 225 125
rect 191 91 225 119
rect 191 51 225 53
rect 191 19 225 51
rect 191 -51 225 -19
rect 191 -53 225 -51
rect 191 -119 225 -91
rect 191 -125 225 -119
rect 191 -187 225 -163
rect 191 -197 225 -187
rect -157 -297 -155 -263
rect -155 -297 -123 -263
rect -85 -297 -53 -263
rect -53 -297 -51 -263
rect 51 -297 53 -263
rect 53 -297 85 -263
rect 123 -297 155 -263
rect 155 -297 157 -263
<< metal1 >>
rect -175 297 -33 303
rect -175 263 -157 297
rect -123 263 -85 297
rect -51 263 -33 297
rect -175 257 -33 263
rect 33 297 175 303
rect 33 263 51 297
rect 85 263 123 297
rect 157 263 175 297
rect 33 257 175 263
rect -231 197 -185 225
rect -231 163 -225 197
rect -191 163 -185 197
rect -231 125 -185 163
rect -231 91 -225 125
rect -191 91 -185 125
rect -231 53 -185 91
rect -231 19 -225 53
rect -191 19 -185 53
rect -231 -19 -185 19
rect -231 -53 -225 -19
rect -191 -53 -185 -19
rect -231 -91 -185 -53
rect -231 -125 -225 -91
rect -191 -125 -185 -91
rect -231 -163 -185 -125
rect -231 -197 -225 -163
rect -191 -197 -185 -163
rect -231 -225 -185 -197
rect -23 197 23 225
rect -23 163 -17 197
rect 17 163 23 197
rect -23 125 23 163
rect -23 91 -17 125
rect 17 91 23 125
rect -23 53 23 91
rect -23 19 -17 53
rect 17 19 23 53
rect -23 -19 23 19
rect -23 -53 -17 -19
rect 17 -53 23 -19
rect -23 -91 23 -53
rect -23 -125 -17 -91
rect 17 -125 23 -91
rect -23 -163 23 -125
rect -23 -197 -17 -163
rect 17 -197 23 -163
rect -23 -225 23 -197
rect 185 197 231 225
rect 185 163 191 197
rect 225 163 231 197
rect 185 125 231 163
rect 185 91 191 125
rect 225 91 231 125
rect 185 53 231 91
rect 185 19 191 53
rect 225 19 231 53
rect 185 -19 231 19
rect 185 -53 191 -19
rect 225 -53 231 -19
rect 185 -91 231 -53
rect 185 -125 191 -91
rect 225 -125 231 -91
rect 185 -163 231 -125
rect 185 -197 191 -163
rect 225 -197 231 -163
rect 185 -225 231 -197
rect -175 -263 -33 -257
rect -175 -297 -157 -263
rect -123 -297 -85 -263
rect -51 -297 -33 -263
rect -175 -303 -33 -297
rect 33 -263 175 -257
rect 33 -297 51 -263
rect 85 -297 123 -263
rect 157 -297 175 -263
rect 33 -303 175 -297
<< properties >>
string FIXED_BBOX -322 -382 322 382
<< end >>
