magic
tech sky130A
magscale 1 2
timestamp 1712816020
<< locali >>
rect 4772 2312 4818 2324
rect 4772 2278 4778 2312
rect 4812 2278 4818 2312
rect 7830 2320 7888 2332
rect 4772 2240 4818 2278
rect 4772 2206 4778 2240
rect 4812 2206 4818 2240
rect 4772 2194 4818 2206
rect 5798 2299 5836 2308
rect 5798 2265 5800 2299
rect 5834 2265 5836 2299
rect 5798 2227 5836 2265
rect 5798 2193 5800 2227
rect 5834 2193 5836 2227
rect 5798 2184 5836 2193
rect 6810 2293 6868 2310
rect 6810 2259 6822 2293
rect 6856 2259 6868 2293
rect 6810 2221 6868 2259
rect 6810 2187 6822 2221
rect 6856 2187 6868 2221
rect 7830 2286 7842 2320
rect 7876 2286 7888 2320
rect 7830 2248 7888 2286
rect 7830 2214 7842 2248
rect 7876 2214 7888 2248
rect 7830 2202 7888 2214
rect 6810 2170 6868 2187
rect 5910 983 5962 984
rect 5910 949 5919 983
rect 5953 949 5962 983
rect 5910 911 5962 949
rect 5910 877 5919 911
rect 5953 877 5962 911
rect 7116 964 7170 988
rect 7116 930 7126 964
rect 7160 930 7170 964
rect 7116 906 7170 930
rect 8336 970 8376 996
rect 8336 936 8339 970
rect 8373 936 8376 970
rect 8336 910 8376 936
rect 9208 976 9272 1002
rect 9208 942 9223 976
rect 9257 942 9272 976
rect 9208 916 9272 942
rect 5910 876 5962 877
rect 4774 624 4830 648
rect 4774 590 4785 624
rect 4819 590 4830 624
rect 4774 552 4830 590
rect 4774 518 4785 552
rect 4819 518 4830 552
rect 4774 494 4830 518
rect 8184 -256 8222 -250
rect 6964 -267 7000 -264
rect 5758 -309 5812 -276
rect 5758 -343 5768 -309
rect 5802 -343 5812 -309
rect 5758 -376 5812 -343
rect 6964 -301 6965 -267
rect 6999 -301 7000 -267
rect 6964 -339 7000 -301
rect 6964 -373 6965 -339
rect 6999 -373 7000 -339
rect 8184 -290 8186 -256
rect 8220 -290 8222 -256
rect 8184 -328 8222 -290
rect 8184 -362 8186 -328
rect 8220 -362 8222 -328
rect 8184 -368 8222 -362
rect 9132 -317 9186 -282
rect 9132 -351 9142 -317
rect 9176 -351 9186 -317
rect 6964 -376 7000 -373
rect 9132 -386 9186 -351
rect 5746 -1418 5800 -1406
rect 5746 -1452 5756 -1418
rect 5790 -1452 5800 -1418
rect 5746 -1490 5800 -1452
rect 5746 -1524 5756 -1490
rect 5790 -1524 5800 -1490
rect 5746 -1536 5800 -1524
rect 6970 -1407 7030 -1376
rect 6970 -1441 6983 -1407
rect 7017 -1441 7030 -1407
rect 6970 -1479 7030 -1441
rect 6970 -1513 6983 -1479
rect 7017 -1513 7030 -1479
rect 6970 -1544 7030 -1513
rect 8176 -1411 8236 -1380
rect 8176 -1445 8189 -1411
rect 8223 -1445 8236 -1411
rect 8176 -1483 8236 -1445
rect 8176 -1517 8189 -1483
rect 8223 -1517 8236 -1483
rect 8176 -1548 8236 -1517
<< viali >>
rect 4778 2278 4812 2312
rect 4778 2206 4812 2240
rect 5800 2265 5834 2299
rect 5800 2193 5834 2227
rect 6822 2259 6856 2293
rect 6822 2187 6856 2221
rect 7842 2286 7876 2320
rect 7842 2214 7876 2248
rect 5919 949 5953 983
rect 5919 877 5953 911
rect 7126 930 7160 964
rect 8339 936 8373 970
rect 9223 942 9257 976
rect 4785 590 4819 624
rect 4785 518 4819 552
rect 5768 -343 5802 -309
rect 6965 -301 6999 -267
rect 6965 -373 6999 -339
rect 8186 -290 8220 -256
rect 8186 -362 8220 -328
rect 9142 -351 9176 -317
rect 5756 -1452 5790 -1418
rect 5756 -1524 5790 -1490
rect 6983 -1441 7017 -1407
rect 6983 -1513 7017 -1479
rect 8189 -1445 8223 -1411
rect 8189 -1517 8223 -1483
<< metal1 >>
rect 5948 2734 6148 2934
rect 5964 2706 6120 2734
rect 5956 2690 6126 2706
rect 5956 2574 5983 2690
rect 6099 2574 6126 2690
rect 5956 2558 6126 2574
rect 4008 2438 4080 2440
rect 4008 2364 7716 2438
rect 4008 1652 4080 2364
rect 4204 2327 4276 2332
rect 4204 2275 4214 2327
rect 4266 2275 4276 2327
rect 4204 2263 4276 2275
rect 4204 2211 4214 2263
rect 4266 2211 4276 2263
rect 4204 2206 4276 2211
rect 4432 2208 4488 2364
rect 4642 2327 4714 2332
rect 4642 2275 4652 2327
rect 4704 2275 4714 2327
rect 4642 2263 4714 2275
rect 4642 2211 4652 2263
rect 4704 2211 4714 2263
rect 4642 2206 4714 2211
rect 4754 2317 4836 2336
rect 7824 2332 7894 2344
rect 5670 2321 5742 2326
rect 4754 2265 4769 2317
rect 4821 2265 4836 2317
rect 4754 2253 4836 2265
rect 4754 2201 4769 2253
rect 4821 2201 4836 2253
rect 4754 2182 4836 2201
rect 5232 2313 5304 2318
rect 5232 2261 5242 2313
rect 5294 2261 5304 2313
rect 5232 2249 5304 2261
rect 5232 2197 5242 2249
rect 5294 2197 5304 2249
rect 5670 2269 5680 2321
rect 5732 2269 5742 2321
rect 5670 2257 5742 2269
rect 5670 2205 5680 2257
rect 5732 2205 5742 2257
rect 5670 2200 5742 2205
rect 5782 2309 5862 2330
rect 5782 2257 5796 2309
rect 5848 2257 5862 2309
rect 5782 2245 5862 2257
rect 5232 2192 5304 2197
rect 5782 2193 5796 2245
rect 5848 2193 5862 2245
rect 5782 2172 5862 2193
rect 6242 2306 6320 2318
rect 6242 2254 6255 2306
rect 6307 2254 6320 2306
rect 6242 2242 6320 2254
rect 6242 2190 6255 2242
rect 6307 2190 6320 2242
rect 6242 2178 6320 2190
rect 6694 2314 6772 2326
rect 7820 2325 7898 2332
rect 6694 2262 6707 2314
rect 6759 2262 6772 2314
rect 6804 2310 6874 2322
rect 7268 2319 7340 2324
rect 6694 2250 6772 2262
rect 6694 2198 6707 2250
rect 6759 2198 6772 2250
rect 6694 2186 6772 2198
rect 6800 2298 6878 2310
rect 6800 2246 6813 2298
rect 6865 2246 6878 2298
rect 6800 2234 6878 2246
rect 6800 2182 6813 2234
rect 6865 2182 6878 2234
rect 7268 2267 7278 2319
rect 7330 2267 7340 2319
rect 7268 2255 7340 2267
rect 7268 2203 7278 2255
rect 7330 2203 7340 2255
rect 7268 2198 7340 2203
rect 7712 2315 7784 2320
rect 7712 2263 7722 2315
rect 7774 2263 7784 2315
rect 7712 2251 7784 2263
rect 7712 2199 7722 2251
rect 7774 2199 7784 2251
rect 7820 2273 7833 2325
rect 7885 2273 7898 2325
rect 7820 2261 7898 2273
rect 7820 2209 7833 2261
rect 7885 2209 7898 2261
rect 7820 2202 7898 2209
rect 7712 2194 7784 2199
rect 7824 2190 7894 2202
rect 6800 2170 6878 2182
rect 6804 2158 6874 2170
rect 4422 1812 4500 1824
rect 4422 1760 4435 1812
rect 4487 1760 4500 1812
rect 4422 1748 4500 1760
rect 4422 1696 4435 1748
rect 4487 1696 4500 1748
rect 4422 1684 4500 1696
rect 5446 1823 5526 1844
rect 5446 1771 5460 1823
rect 5512 1771 5526 1823
rect 5446 1759 5526 1771
rect 5446 1707 5460 1759
rect 5512 1707 5526 1759
rect 5446 1686 5526 1707
rect 6472 1813 6548 1818
rect 6472 1761 6484 1813
rect 6536 1761 6548 1813
rect 6472 1749 6548 1761
rect 6472 1697 6484 1749
rect 6536 1697 6548 1749
rect 6472 1692 6548 1697
rect 7494 1775 7572 1804
rect 7494 1723 7507 1775
rect 7559 1723 7572 1775
rect 7494 1694 7572 1723
rect 4008 1578 7722 1652
rect 4008 1576 4080 1578
rect 8294 1447 8396 1460
rect 7094 1442 7200 1444
rect 8294 1442 8319 1447
rect 5878 1438 8319 1442
rect 5878 1436 7121 1438
rect 5878 1384 5905 1436
rect 5957 1386 7121 1436
rect 7173 1395 8319 1438
rect 8371 1395 8396 1447
rect 7173 1386 8396 1395
rect 5957 1384 8396 1386
rect 5878 1382 8396 1384
rect 5878 1378 8366 1382
rect 4954 1334 5128 1338
rect 4954 1332 6196 1334
rect 8630 1332 8696 1336
rect 4954 1330 7374 1332
rect 8516 1330 8696 1332
rect 4954 1270 8696 1330
rect 4026 1222 4108 1224
rect 4026 1156 4664 1222
rect 4026 778 4108 1156
rect 4432 1093 4504 1124
rect 4432 1041 4442 1093
rect 4494 1041 4504 1093
rect 4432 1010 4504 1041
rect 4958 1082 5026 1270
rect 5090 1268 8696 1270
rect 5090 1266 8524 1268
rect 6196 1264 8524 1266
rect 7366 1260 8524 1264
rect 8630 1098 8696 1268
rect 8630 1096 9008 1098
rect 7440 1082 8208 1084
rect 4958 1028 5792 1082
rect 6162 1028 6996 1082
rect 7374 1030 8208 1082
rect 8628 1038 9008 1096
rect 4958 1012 5026 1028
rect 3508 580 4108 778
rect 4768 648 4836 660
rect 3508 578 3708 580
rect 3760 -1030 3952 580
rect 4026 450 4108 580
rect 4208 617 4298 630
rect 4208 565 4227 617
rect 4279 565 4298 617
rect 4208 553 4298 565
rect 4208 501 4227 553
rect 4279 501 4298 553
rect 4208 488 4298 501
rect 4646 629 4736 642
rect 4646 577 4665 629
rect 4717 577 4736 629
rect 4646 565 4736 577
rect 4646 513 4665 565
rect 4717 513 4736 565
rect 4646 500 4736 513
rect 4764 629 4840 648
rect 4764 577 4776 629
rect 4828 577 4840 629
rect 4764 565 4840 577
rect 4764 513 4776 565
rect 4828 513 4840 565
rect 4764 494 4840 513
rect 4958 550 5024 1012
rect 5160 954 5232 982
rect 5160 902 5170 954
rect 5222 902 5232 954
rect 5160 874 5232 902
rect 5572 960 5644 988
rect 5904 984 5968 996
rect 5572 908 5582 960
rect 5634 908 5644 960
rect 5572 880 5644 908
rect 5900 983 5972 984
rect 5900 956 5919 983
rect 5953 956 5972 983
rect 5900 904 5910 956
rect 5962 904 5972 956
rect 5900 877 5919 904
rect 5953 877 5972 904
rect 5900 876 5972 877
rect 5904 864 5968 876
rect 5370 668 5442 692
rect 5370 616 5380 668
rect 5432 616 5442 668
rect 5370 592 5442 616
rect 5786 668 5858 692
rect 5786 616 5796 668
rect 5848 616 5858 668
rect 5786 592 5858 616
rect 6162 550 6228 1028
rect 6370 975 6444 990
rect 6370 923 6381 975
rect 6433 923 6444 975
rect 6370 908 6444 923
rect 6784 977 6858 992
rect 7110 988 7176 1000
rect 6784 925 6795 977
rect 6847 925 6858 977
rect 6784 910 6858 925
rect 7106 973 7180 988
rect 7106 921 7117 973
rect 7169 921 7180 973
rect 7106 906 7180 921
rect 7110 894 7176 906
rect 6578 660 6654 680
rect 6578 608 6590 660
rect 6642 608 6654 660
rect 6578 588 6654 608
rect 6994 668 7070 688
rect 6994 616 7006 668
rect 7058 616 7070 668
rect 6994 596 7070 616
rect 7374 552 7440 1030
rect 8330 998 8382 1008
rect 7574 971 7658 988
rect 7574 919 7590 971
rect 7642 919 7658 971
rect 7574 902 7658 919
rect 7994 977 8078 994
rect 7994 925 8010 977
rect 8062 925 8078 977
rect 7994 908 8078 925
rect 8322 977 8394 998
rect 8322 925 8332 977
rect 8384 925 8394 977
rect 8322 904 8394 925
rect 8330 898 8382 904
rect 7784 664 7864 682
rect 7784 612 7798 664
rect 7850 612 7864 664
rect 7784 594 7864 612
rect 8208 658 8288 676
rect 8208 606 8222 658
rect 8274 606 8288 658
rect 8628 650 8696 1038
rect 8792 987 8876 1004
rect 9202 1002 9278 1014
rect 8792 935 8808 987
rect 8860 935 8876 987
rect 8792 918 8876 935
rect 8982 985 9066 1002
rect 8982 933 8998 985
rect 9050 933 9066 985
rect 8982 916 9066 933
rect 9198 985 9282 1002
rect 9198 933 9214 985
rect 9266 933 9282 985
rect 9198 916 9282 933
rect 9202 904 9278 916
rect 8208 588 8288 606
rect 8626 570 8696 650
rect 8892 682 8964 698
rect 8892 630 8902 682
rect 8954 630 8964 682
rect 8892 614 8964 630
rect 9086 688 9158 704
rect 9086 636 9096 688
rect 9148 636 9158 688
rect 9086 620 9158 636
rect 4958 496 5792 550
rect 6162 496 6996 550
rect 7374 498 8208 552
rect 8626 510 9100 570
rect 8626 506 8696 510
rect 4768 482 4836 494
rect 4026 384 4654 450
rect 4026 382 4108 384
rect 4958 152 5024 496
rect 6162 362 6228 496
rect 6148 358 6236 362
rect 6148 306 6166 358
rect 6218 306 6236 358
rect 7374 354 7440 498
rect 8626 366 8694 506
rect 8898 392 8998 396
rect 9378 392 9578 434
rect 8898 374 9578 392
rect 6632 352 7440 354
rect 6148 302 6236 306
rect 6620 350 7440 352
rect 6162 152 6228 302
rect 6620 298 6636 350
rect 6688 298 7440 350
rect 6620 296 6704 298
rect 7374 154 7440 298
rect 8616 354 8702 366
rect 8616 302 8633 354
rect 8685 302 8702 354
rect 8616 290 8702 302
rect 8898 322 8922 374
rect 8974 322 9578 374
rect 8898 300 9578 322
rect 8916 292 9578 300
rect 4958 98 5636 152
rect 6162 98 6840 152
rect 7374 100 8052 154
rect 8626 138 8694 290
rect 9378 234 9578 292
rect 4958 -412 5024 98
rect 5422 47 5496 66
rect 5422 -5 5433 47
rect 5485 -5 5496 47
rect 5422 -24 5496 -5
rect 5216 -296 5290 -272
rect 5216 -348 5227 -296
rect 5279 -348 5290 -296
rect 5216 -372 5290 -348
rect 5630 -294 5704 -270
rect 5752 -274 5818 -264
rect 5630 -346 5641 -294
rect 5693 -346 5704 -294
rect 5630 -370 5704 -346
rect 5748 -300 5992 -274
rect 5748 -352 5759 -300
rect 5811 -352 5992 -300
rect 5748 -384 5992 -352
rect 5752 -388 5818 -384
rect 4958 -466 5638 -412
rect 4412 -598 4538 -594
rect 5862 -598 5990 -384
rect 6162 -414 6228 98
rect 6622 47 6700 66
rect 6622 -5 6635 47
rect 6687 -5 6700 47
rect 6622 -24 6700 -5
rect 6958 -264 7006 -252
rect 6944 -265 7020 -264
rect 6414 -302 6488 -278
rect 6414 -354 6425 -302
rect 6477 -354 6488 -302
rect 6414 -378 6488 -354
rect 6830 -295 6908 -266
rect 6830 -347 6843 -295
rect 6895 -347 6908 -295
rect 6830 -376 6908 -347
rect 6944 -317 6956 -265
rect 7008 -270 7020 -265
rect 7058 -270 7154 -268
rect 7008 -317 7154 -270
rect 6944 -329 7154 -317
rect 6944 -381 6956 -329
rect 7008 -380 7154 -329
rect 7008 -381 7020 -380
rect 6944 -382 7020 -381
rect 6958 -388 7006 -382
rect 6162 -468 6842 -414
rect 4412 -602 5990 -598
rect 7058 -602 7154 -380
rect 7374 -410 7440 100
rect 8626 90 9028 138
rect 7842 36 7914 66
rect 7842 -16 7852 36
rect 7904 -16 7914 36
rect 7842 -46 7914 -16
rect 8178 -242 8228 -238
rect 8308 -242 8392 -240
rect 8164 -251 8392 -242
rect 7632 -292 7704 -262
rect 7632 -344 7642 -292
rect 7694 -344 7704 -292
rect 7632 -374 7704 -344
rect 8052 -286 8124 -256
rect 8052 -338 8062 -286
rect 8114 -338 8124 -286
rect 8052 -368 8124 -338
rect 8164 -303 8175 -251
rect 8227 -303 8392 -251
rect 8164 -315 8392 -303
rect 8164 -367 8175 -315
rect 8227 -367 8392 -315
rect 8164 -372 8392 -367
rect 8164 -376 8238 -372
rect 8178 -380 8228 -376
rect 7374 -464 8054 -410
rect 8308 -602 8392 -372
rect 8626 -424 8694 90
rect 8726 86 9028 90
rect 8912 20 8984 50
rect 8912 -32 8922 20
rect 8974 -32 8984 20
rect 8912 -62 8984 -32
rect 9126 -282 9192 -270
rect 8820 -312 8894 -286
rect 8820 -364 8831 -312
rect 8883 -364 8894 -312
rect 8820 -390 8894 -364
rect 9012 -314 9086 -288
rect 9012 -366 9023 -314
rect 9075 -366 9086 -314
rect 9012 -392 9086 -366
rect 9122 -308 9196 -282
rect 9122 -360 9133 -308
rect 9185 -360 9196 -308
rect 9122 -386 9196 -360
rect 9126 -398 9192 -386
rect 8626 -484 8932 -424
rect 4412 -606 8392 -602
rect 4412 -658 4449 -606
rect 4501 -658 8392 -606
rect 4412 -668 8392 -658
rect 4412 -670 5990 -668
rect 4904 -786 5004 -784
rect 4904 -872 8078 -786
rect 4904 -1030 5004 -872
rect 3760 -1220 5004 -1030
rect 5390 -949 5468 -918
rect 5390 -1001 5403 -949
rect 5455 -1001 5468 -949
rect 5390 -1032 5468 -1001
rect 6614 -932 6696 -902
rect 6614 -984 6629 -932
rect 6681 -984 6696 -932
rect 6614 -1014 6696 -984
rect 7838 -934 7914 -908
rect 7838 -986 7850 -934
rect 7902 -986 7914 -934
rect 7838 -1012 7914 -986
rect 4904 -1584 5004 -1220
rect 5740 -1406 5806 -1394
rect 5624 -1413 5698 -1406
rect 5184 -1425 5258 -1418
rect 5184 -1477 5195 -1425
rect 5247 -1477 5258 -1425
rect 5184 -1489 5258 -1477
rect 5184 -1541 5195 -1489
rect 5247 -1541 5258 -1489
rect 5624 -1465 5635 -1413
rect 5687 -1465 5698 -1413
rect 5624 -1477 5698 -1465
rect 5624 -1529 5635 -1477
rect 5687 -1529 5698 -1477
rect 5624 -1536 5698 -1529
rect 5736 -1413 5810 -1406
rect 5736 -1465 5747 -1413
rect 5799 -1465 5810 -1413
rect 5736 -1477 5810 -1465
rect 5736 -1529 5747 -1477
rect 5799 -1529 5810 -1477
rect 5736 -1536 5810 -1529
rect 6400 -1408 6480 -1382
rect 6400 -1460 6414 -1408
rect 6466 -1460 6480 -1408
rect 6400 -1472 6480 -1460
rect 6400 -1524 6414 -1472
rect 6466 -1524 6480 -1472
rect 5184 -1548 5258 -1541
rect 5740 -1548 5806 -1536
rect 6400 -1550 6480 -1524
rect 6842 -1396 6922 -1370
rect 6964 -1376 7036 -1364
rect 6842 -1448 6856 -1396
rect 6908 -1448 6922 -1396
rect 6842 -1460 6922 -1448
rect 6842 -1512 6856 -1460
rect 6908 -1512 6922 -1460
rect 6842 -1538 6922 -1512
rect 6960 -1402 7040 -1376
rect 6960 -1454 6974 -1402
rect 7026 -1454 7040 -1402
rect 6960 -1466 7040 -1454
rect 6960 -1518 6974 -1466
rect 7026 -1518 7040 -1466
rect 6960 -1544 7040 -1518
rect 7622 -1402 7702 -1376
rect 7622 -1454 7636 -1402
rect 7688 -1454 7702 -1402
rect 7622 -1466 7702 -1454
rect 7622 -1518 7636 -1466
rect 7688 -1518 7702 -1466
rect 7622 -1544 7702 -1518
rect 8054 -1404 8134 -1378
rect 8170 -1380 8242 -1368
rect 8054 -1456 8068 -1404
rect 8120 -1456 8134 -1404
rect 8054 -1468 8134 -1456
rect 8054 -1520 8068 -1468
rect 8120 -1520 8134 -1468
rect 6964 -1556 7036 -1544
rect 8054 -1546 8134 -1520
rect 8166 -1406 8246 -1380
rect 8166 -1458 8180 -1406
rect 8232 -1458 8246 -1406
rect 8166 -1470 8246 -1458
rect 8166 -1522 8180 -1470
rect 8232 -1522 8246 -1470
rect 8166 -1548 8246 -1522
rect 8170 -1560 8242 -1548
rect 4904 -1662 8074 -1584
rect 4910 -1670 8074 -1662
rect 7090 -1823 7312 -1804
rect 7090 -1939 7111 -1823
rect 7291 -1939 7312 -1823
rect 7090 -1958 7312 -1939
rect 7098 -2212 7298 -1958
<< via1 >>
rect 5983 2574 6099 2690
rect 4214 2275 4266 2327
rect 4214 2211 4266 2263
rect 4652 2275 4704 2327
rect 4652 2211 4704 2263
rect 4769 2312 4821 2317
rect 4769 2278 4778 2312
rect 4778 2278 4812 2312
rect 4812 2278 4821 2312
rect 4769 2265 4821 2278
rect 4769 2240 4821 2253
rect 4769 2206 4778 2240
rect 4778 2206 4812 2240
rect 4812 2206 4821 2240
rect 4769 2201 4821 2206
rect 5242 2261 5294 2313
rect 5242 2197 5294 2249
rect 5680 2269 5732 2321
rect 5680 2205 5732 2257
rect 5796 2299 5848 2309
rect 5796 2265 5800 2299
rect 5800 2265 5834 2299
rect 5834 2265 5848 2299
rect 5796 2257 5848 2265
rect 5796 2227 5848 2245
rect 5796 2193 5800 2227
rect 5800 2193 5834 2227
rect 5834 2193 5848 2227
rect 6255 2254 6307 2306
rect 6255 2190 6307 2242
rect 6707 2262 6759 2314
rect 6707 2198 6759 2250
rect 6813 2293 6865 2298
rect 6813 2259 6822 2293
rect 6822 2259 6856 2293
rect 6856 2259 6865 2293
rect 6813 2246 6865 2259
rect 6813 2221 6865 2234
rect 6813 2187 6822 2221
rect 6822 2187 6856 2221
rect 6856 2187 6865 2221
rect 6813 2182 6865 2187
rect 7278 2267 7330 2319
rect 7278 2203 7330 2255
rect 7722 2263 7774 2315
rect 7722 2199 7774 2251
rect 7833 2320 7885 2325
rect 7833 2286 7842 2320
rect 7842 2286 7876 2320
rect 7876 2286 7885 2320
rect 7833 2273 7885 2286
rect 7833 2248 7885 2261
rect 7833 2214 7842 2248
rect 7842 2214 7876 2248
rect 7876 2214 7885 2248
rect 7833 2209 7885 2214
rect 4435 1760 4487 1812
rect 4435 1696 4487 1748
rect 5460 1771 5512 1823
rect 5460 1707 5512 1759
rect 6484 1761 6536 1813
rect 6484 1697 6536 1749
rect 7507 1723 7559 1775
rect 5905 1384 5957 1436
rect 7121 1386 7173 1438
rect 8319 1395 8371 1447
rect 4442 1041 4494 1093
rect 4227 565 4279 617
rect 4227 501 4279 553
rect 4665 577 4717 629
rect 4665 513 4717 565
rect 4776 624 4828 629
rect 4776 590 4785 624
rect 4785 590 4819 624
rect 4819 590 4828 624
rect 4776 577 4828 590
rect 4776 552 4828 565
rect 4776 518 4785 552
rect 4785 518 4819 552
rect 4819 518 4828 552
rect 4776 513 4828 518
rect 5170 902 5222 954
rect 5582 908 5634 960
rect 5910 949 5919 956
rect 5919 949 5953 956
rect 5953 949 5962 956
rect 5910 911 5962 949
rect 5910 904 5919 911
rect 5919 904 5953 911
rect 5953 904 5962 911
rect 5380 616 5432 668
rect 5796 616 5848 668
rect 6381 923 6433 975
rect 6795 925 6847 977
rect 7117 964 7169 973
rect 7117 930 7126 964
rect 7126 930 7160 964
rect 7160 930 7169 964
rect 7117 921 7169 930
rect 6590 608 6642 660
rect 7006 616 7058 668
rect 7590 919 7642 971
rect 8010 925 8062 977
rect 8332 970 8384 977
rect 8332 936 8339 970
rect 8339 936 8373 970
rect 8373 936 8384 970
rect 8332 925 8384 936
rect 7798 612 7850 664
rect 8222 606 8274 658
rect 8808 935 8860 987
rect 8998 933 9050 985
rect 9214 976 9266 985
rect 9214 942 9223 976
rect 9223 942 9257 976
rect 9257 942 9266 976
rect 9214 933 9266 942
rect 8902 630 8954 682
rect 9096 636 9148 688
rect 6166 306 6218 358
rect 6636 298 6688 350
rect 8633 302 8685 354
rect 8922 322 8974 374
rect 5433 -5 5485 47
rect 5227 -348 5279 -296
rect 5641 -346 5693 -294
rect 5759 -309 5811 -300
rect 5759 -343 5768 -309
rect 5768 -343 5802 -309
rect 5802 -343 5811 -309
rect 5759 -352 5811 -343
rect 6635 -5 6687 47
rect 6425 -354 6477 -302
rect 6843 -347 6895 -295
rect 6956 -267 7008 -265
rect 6956 -301 6965 -267
rect 6965 -301 6999 -267
rect 6999 -301 7008 -267
rect 6956 -317 7008 -301
rect 6956 -339 7008 -329
rect 6956 -373 6965 -339
rect 6965 -373 6999 -339
rect 6999 -373 7008 -339
rect 6956 -381 7008 -373
rect 7852 -16 7904 36
rect 7642 -344 7694 -292
rect 8062 -338 8114 -286
rect 8175 -256 8227 -251
rect 8175 -290 8186 -256
rect 8186 -290 8220 -256
rect 8220 -290 8227 -256
rect 8175 -303 8227 -290
rect 8175 -328 8227 -315
rect 8175 -362 8186 -328
rect 8186 -362 8220 -328
rect 8220 -362 8227 -328
rect 8175 -367 8227 -362
rect 8922 -32 8974 20
rect 8831 -364 8883 -312
rect 9023 -366 9075 -314
rect 9133 -317 9185 -308
rect 9133 -351 9142 -317
rect 9142 -351 9176 -317
rect 9176 -351 9185 -317
rect 9133 -360 9185 -351
rect 4449 -658 4501 -606
rect 5403 -1001 5455 -949
rect 6629 -984 6681 -932
rect 7850 -986 7902 -934
rect 5195 -1477 5247 -1425
rect 5195 -1541 5247 -1489
rect 5635 -1465 5687 -1413
rect 5635 -1529 5687 -1477
rect 5747 -1418 5799 -1413
rect 5747 -1452 5756 -1418
rect 5756 -1452 5790 -1418
rect 5790 -1452 5799 -1418
rect 5747 -1465 5799 -1452
rect 5747 -1490 5799 -1477
rect 5747 -1524 5756 -1490
rect 5756 -1524 5790 -1490
rect 5790 -1524 5799 -1490
rect 5747 -1529 5799 -1524
rect 6414 -1460 6466 -1408
rect 6414 -1524 6466 -1472
rect 6856 -1448 6908 -1396
rect 6856 -1512 6908 -1460
rect 6974 -1407 7026 -1402
rect 6974 -1441 6983 -1407
rect 6983 -1441 7017 -1407
rect 7017 -1441 7026 -1407
rect 6974 -1454 7026 -1441
rect 6974 -1479 7026 -1466
rect 6974 -1513 6983 -1479
rect 6983 -1513 7017 -1479
rect 7017 -1513 7026 -1479
rect 6974 -1518 7026 -1513
rect 7636 -1454 7688 -1402
rect 7636 -1518 7688 -1466
rect 8068 -1456 8120 -1404
rect 8068 -1520 8120 -1468
rect 8180 -1411 8232 -1406
rect 8180 -1445 8189 -1411
rect 8189 -1445 8223 -1411
rect 8223 -1445 8232 -1411
rect 8180 -1458 8232 -1445
rect 8180 -1483 8232 -1470
rect 8180 -1517 8189 -1483
rect 8189 -1517 8223 -1483
rect 8223 -1517 8232 -1483
rect 8180 -1522 8232 -1517
rect 7111 -1939 7291 -1823
<< metal2 >>
rect 8862 2722 9006 2726
rect 5984 2716 9006 2722
rect 5966 2690 9006 2716
rect 5966 2642 5983 2690
rect 5964 2574 5983 2642
rect 6099 2574 9006 2690
rect 5964 2570 9006 2574
rect 4214 2332 4266 2342
rect 4652 2332 4704 2342
rect 4764 2332 4826 2346
rect 5680 2332 5732 2336
rect 5792 2332 5852 2340
rect 5964 2332 6116 2570
rect 6704 2332 6762 2336
rect 7278 2332 7330 2334
rect 7830 2332 7888 2342
rect 4196 2327 7888 2332
rect 4196 2275 4214 2327
rect 4266 2275 4652 2327
rect 4704 2325 7888 2327
rect 4704 2321 7833 2325
rect 4704 2317 5680 2321
rect 4704 2275 4769 2317
rect 4196 2265 4769 2275
rect 4821 2313 5680 2317
rect 4821 2265 5242 2313
rect 4196 2263 5242 2265
rect 4196 2211 4214 2263
rect 4266 2211 4652 2263
rect 4704 2261 5242 2263
rect 5294 2269 5680 2313
rect 5732 2319 7833 2321
rect 5732 2314 7278 2319
rect 5732 2309 6707 2314
rect 5732 2269 5796 2309
rect 5294 2261 5796 2269
rect 4704 2257 5796 2261
rect 5848 2306 6707 2309
rect 5848 2257 6255 2306
rect 4704 2253 5680 2257
rect 4704 2211 4769 2253
rect 4196 2206 4769 2211
rect 4214 2196 4266 2206
rect 4652 2196 4704 2206
rect 4764 2201 4769 2206
rect 4821 2249 5680 2253
rect 4821 2206 5242 2249
rect 4821 2201 4826 2206
rect 4764 2172 4826 2201
rect 5294 2206 5680 2249
rect 5242 2182 5294 2197
rect 5732 2254 6255 2257
rect 6307 2262 6707 2306
rect 6759 2298 7278 2314
rect 6759 2262 6813 2298
rect 6307 2254 6813 2262
rect 5732 2250 6813 2254
rect 5732 2245 6707 2250
rect 5732 2206 5796 2245
rect 5680 2190 5732 2205
rect 5792 2193 5796 2206
rect 5848 2242 6707 2245
rect 5848 2206 6255 2242
rect 5848 2193 5852 2206
rect 5792 2162 5852 2193
rect 6252 2190 6255 2206
rect 6307 2206 6707 2242
rect 6307 2190 6310 2206
rect 6252 2168 6310 2190
rect 6704 2198 6707 2206
rect 6759 2246 6813 2250
rect 6865 2267 7278 2298
rect 7330 2315 7833 2319
rect 7330 2267 7722 2315
rect 6865 2263 7722 2267
rect 7774 2273 7833 2315
rect 7885 2273 7888 2325
rect 7774 2263 7888 2273
rect 6865 2261 7888 2263
rect 6865 2255 7833 2261
rect 6865 2246 7278 2255
rect 6759 2234 7278 2246
rect 6759 2206 6813 2234
rect 6759 2198 6762 2206
rect 6704 2176 6762 2198
rect 6810 2182 6813 2206
rect 6865 2206 7278 2234
rect 6865 2182 6868 2206
rect 7330 2251 7833 2255
rect 7330 2206 7722 2251
rect 7278 2188 7330 2203
rect 7774 2209 7833 2251
rect 7885 2209 7888 2261
rect 7774 2206 7888 2209
rect 7722 2184 7774 2199
rect 7830 2192 7888 2206
rect 6810 2160 6868 2182
rect 5456 1850 5516 1854
rect 4432 1824 4490 1834
rect 4432 1812 4498 1824
rect 4432 1760 4435 1812
rect 4487 1760 4498 1812
rect 4432 1748 4498 1760
rect 4432 1696 4435 1748
rect 4487 1696 4498 1748
rect 4432 1093 4498 1696
rect 4432 1041 4442 1093
rect 4494 1041 4498 1093
rect 4432 1010 4498 1041
rect 5434 1823 5516 1850
rect 6482 1824 6538 1828
rect 5434 1771 5460 1823
rect 5512 1771 5516 1823
rect 5434 1759 5516 1771
rect 5434 1707 5460 1759
rect 5512 1707 5516 1759
rect 5434 1676 5516 1707
rect 6470 1813 6544 1824
rect 6470 1761 6484 1813
rect 6536 1761 6544 1813
rect 6470 1749 6544 1761
rect 6470 1697 6484 1749
rect 6536 1697 6544 1749
rect 7504 1775 7562 1814
rect 7504 1723 7507 1775
rect 7559 1723 7562 1775
rect 7504 1700 7562 1723
rect 4442 1000 4494 1010
rect 5170 976 5222 992
rect 5434 976 5512 1676
rect 5888 1436 5974 1452
rect 5888 1384 5905 1436
rect 5957 1384 5974 1436
rect 5888 1368 5974 1384
rect 5582 976 5634 998
rect 5164 960 5634 976
rect 5164 954 5582 960
rect 5164 902 5170 954
rect 5222 908 5582 954
rect 5222 902 5634 908
rect 5164 872 5634 902
rect 5170 864 5222 872
rect 5582 870 5634 872
rect 5894 956 5972 1368
rect 5894 904 5910 956
rect 5962 904 5972 956
rect 5894 870 5972 904
rect 6380 994 6434 1000
rect 6470 994 6544 1697
rect 7502 1684 7562 1700
rect 7104 1438 7190 1454
rect 7104 1386 7121 1438
rect 7173 1386 7190 1438
rect 7104 1370 7190 1386
rect 6794 994 6848 1002
rect 6380 977 6848 994
rect 6380 975 6795 977
rect 6380 923 6381 975
rect 6433 925 6795 975
rect 6847 925 6848 977
rect 6433 923 6848 925
rect 6380 904 6848 923
rect 6380 898 6434 904
rect 6794 900 6848 904
rect 7106 973 7184 1370
rect 7502 1366 7560 1684
rect 8304 1447 8396 2570
rect 8304 1395 8319 1447
rect 8371 1395 8396 1447
rect 8304 1382 8396 1395
rect 8304 1372 8388 1382
rect 7502 1308 7796 1366
rect 7502 1306 7560 1308
rect 7584 992 7648 998
rect 7724 992 7796 1308
rect 8004 996 8068 1004
rect 8002 992 8068 996
rect 7106 921 7117 973
rect 7169 921 7184 973
rect 7106 896 7184 921
rect 7576 977 8068 992
rect 7576 971 8010 977
rect 7576 919 7590 971
rect 7642 925 8010 971
rect 8062 925 8068 977
rect 7642 919 8068 925
rect 7576 904 8068 919
rect 8310 977 8388 1372
rect 8862 1014 9006 2570
rect 8802 1012 9006 1014
rect 8802 1004 9056 1012
rect 9208 1004 9272 1012
rect 8310 925 8332 977
rect 8384 925 8388 977
rect 8310 908 8388 925
rect 8790 987 9274 1004
rect 8790 935 8808 987
rect 8860 985 9274 987
rect 8860 935 8998 985
rect 8790 933 8998 935
rect 9050 933 9214 985
rect 9266 933 9274 985
rect 8790 918 9274 933
rect 8802 908 8866 918
rect 7584 892 7648 904
rect 8004 898 8068 904
rect 8332 894 8384 908
rect 8992 906 9056 918
rect 9208 906 9272 918
rect 5910 866 5962 870
rect 8902 702 8954 708
rect 9096 702 9148 714
rect 5380 692 5432 702
rect 5796 692 5848 702
rect 5374 668 5848 692
rect 6588 688 6644 690
rect 7004 688 7060 698
rect 4218 634 4288 640
rect 4656 634 4726 652
rect 4774 634 4830 658
rect 4212 629 4832 634
rect 4212 617 4665 629
rect 4212 565 4227 617
rect 4279 577 4665 617
rect 4717 577 4776 629
rect 4828 577 4832 629
rect 5374 616 5380 668
rect 5432 616 5796 668
rect 5374 590 5848 616
rect 5380 582 5496 590
rect 5796 582 5848 590
rect 6586 668 7060 688
rect 6586 660 7006 668
rect 6586 608 6590 660
rect 6642 616 7006 660
rect 7058 616 7060 668
rect 6642 608 7060 616
rect 6586 586 7060 608
rect 7794 680 7854 692
rect 8900 688 9156 702
rect 8218 680 8278 686
rect 7794 664 8278 680
rect 7794 612 7798 664
rect 7850 658 8278 664
rect 7850 612 8222 658
rect 7794 606 8222 612
rect 8274 606 8278 658
rect 8900 682 9096 688
rect 8900 630 8902 682
rect 8954 636 9096 682
rect 9148 636 9156 688
rect 8954 630 9156 636
rect 8900 616 9156 630
rect 7794 600 8278 606
rect 8902 604 8986 616
rect 9096 610 9148 616
rect 4279 565 4832 577
rect 4212 553 4665 565
rect 4212 501 4227 553
rect 4279 513 4665 553
rect 4717 513 4776 565
rect 4828 513 4832 565
rect 4279 501 4832 513
rect 4212 492 4832 501
rect 4218 478 4288 492
rect 4394 -606 4530 492
rect 4656 490 4726 492
rect 4774 484 4830 492
rect 5432 362 5496 582
rect 6588 578 6692 586
rect 7794 584 7914 600
rect 6158 362 6226 372
rect 6632 362 6692 578
rect 7844 364 7914 584
rect 8218 578 8278 600
rect 8914 406 8986 604
rect 8626 364 8692 376
rect 5426 358 6228 362
rect 5426 306 6166 358
rect 6218 306 6228 358
rect 5426 302 6228 306
rect 6630 350 6694 362
rect 5432 47 5496 302
rect 6158 292 6226 302
rect 6630 298 6636 350
rect 6688 298 6694 350
rect 6630 286 6694 298
rect 7844 354 8692 364
rect 7844 302 8633 354
rect 8685 302 8692 354
rect 7844 292 8692 302
rect 7844 290 7914 292
rect 5432 -5 5433 47
rect 5485 -5 5496 47
rect 5432 -24 5496 -5
rect 6632 47 6692 286
rect 6632 -5 6635 47
rect 6687 -5 6692 47
rect 5432 -34 5486 -24
rect 6632 -28 6692 -5
rect 7846 36 7912 290
rect 8626 280 8692 292
rect 8908 374 8988 406
rect 8908 322 8922 374
rect 8974 322 8988 374
rect 8908 290 8988 322
rect 7846 -16 7852 36
rect 7904 -16 7912 36
rect 6632 -34 6690 -28
rect 7846 -46 7912 -16
rect 8914 20 8986 290
rect 8914 -32 8922 20
rect 8974 -32 8986 20
rect 7852 -56 7904 -46
rect 8914 -62 8986 -32
rect 8922 -72 8974 -62
rect 8062 -252 8114 -246
rect 5226 -272 5280 -262
rect 5640 -272 5694 -260
rect 5214 -294 5694 -272
rect 5214 -296 5641 -294
rect 5214 -348 5227 -296
rect 5279 -346 5641 -296
rect 5693 -346 5694 -294
rect 5279 -348 5694 -346
rect 5214 -372 5694 -348
rect 5226 -382 5280 -372
rect 4394 -658 4449 -606
rect 4501 -658 4530 -606
rect 4394 -1806 4530 -658
rect 5396 -924 5462 -372
rect 5640 -380 5694 -372
rect 5758 -272 5812 -266
rect 6424 -270 6478 -268
rect 6840 -270 6898 -256
rect 5758 -300 5824 -272
rect 5758 -352 5759 -300
rect 5811 -352 5824 -300
rect 5758 -372 5824 -352
rect 6422 -295 6898 -270
rect 6422 -302 6843 -295
rect 6422 -354 6425 -302
rect 6477 -347 6843 -302
rect 6895 -347 6898 -295
rect 6477 -354 6898 -347
rect 5758 -386 5812 -372
rect 6422 -378 6898 -354
rect 6424 -388 6478 -378
rect 5396 -949 5458 -924
rect 5396 -1001 5403 -949
rect 5455 -1001 5458 -949
rect 5396 -1036 5458 -1001
rect 6624 -932 6690 -378
rect 6840 -386 6898 -378
rect 6954 -265 7010 -254
rect 6954 -317 6956 -265
rect 7008 -317 7010 -265
rect 6954 -329 7010 -317
rect 6954 -381 6956 -329
rect 7008 -381 7010 -329
rect 7640 -286 8114 -252
rect 7640 -292 8062 -286
rect 7640 -344 7642 -292
rect 7694 -338 8062 -292
rect 7694 -344 8114 -338
rect 7640 -376 8114 -344
rect 6954 -392 7010 -381
rect 7642 -384 7694 -376
rect 6624 -984 6629 -932
rect 6681 -984 6690 -932
rect 6624 -1014 6690 -984
rect 7848 -934 7908 -376
rect 8062 -378 8114 -376
rect 8174 -251 8228 -232
rect 8174 -303 8175 -251
rect 8227 -303 8228 -251
rect 8830 -284 8884 -276
rect 9022 -284 9076 -278
rect 9132 -284 9186 -272
rect 8174 -315 8228 -303
rect 8174 -367 8175 -315
rect 8227 -367 8228 -315
rect 8174 -386 8228 -367
rect 8826 -308 9192 -284
rect 8826 -312 9133 -308
rect 8826 -364 8831 -312
rect 8883 -314 9133 -312
rect 8883 -364 9023 -314
rect 8826 -366 9023 -364
rect 9075 -360 9133 -314
rect 9185 -360 9192 -308
rect 9075 -366 9192 -360
rect 8826 -392 9192 -366
rect 8830 -400 8982 -392
rect 7848 -986 7850 -934
rect 7902 -986 7908 -934
rect 7848 -1012 7908 -986
rect 6624 -1024 6686 -1014
rect 7848 -1022 7904 -1012
rect 5400 -1042 5458 -1036
rect 6410 -1382 6470 -1372
rect 6852 -1382 6912 -1360
rect 6970 -1382 7030 -1366
rect 7632 -1382 7692 -1366
rect 8064 -1382 8124 -1368
rect 8176 -1382 8236 -1370
rect 5184 -1396 8248 -1382
rect 5184 -1408 6856 -1396
rect 5184 -1413 6414 -1408
rect 5184 -1425 5635 -1413
rect 5184 -1477 5195 -1425
rect 5247 -1465 5635 -1425
rect 5687 -1465 5747 -1413
rect 5799 -1460 6414 -1413
rect 6466 -1448 6856 -1408
rect 6908 -1402 8248 -1396
rect 6908 -1448 6974 -1402
rect 6466 -1454 6974 -1448
rect 7026 -1454 7636 -1402
rect 7688 -1404 8248 -1402
rect 7688 -1454 8068 -1404
rect 6466 -1456 8068 -1454
rect 8120 -1406 8248 -1404
rect 8120 -1456 8180 -1406
rect 6466 -1458 8180 -1456
rect 8232 -1458 8248 -1406
rect 6466 -1460 8248 -1458
rect 5799 -1465 6856 -1460
rect 5247 -1472 6856 -1465
rect 5247 -1477 6414 -1472
rect 5184 -1489 5635 -1477
rect 5184 -1541 5195 -1489
rect 5247 -1529 5635 -1489
rect 5687 -1529 5747 -1477
rect 5799 -1524 6414 -1477
rect 6466 -1512 6856 -1472
rect 6908 -1466 8248 -1460
rect 6908 -1512 6974 -1466
rect 6466 -1518 6974 -1512
rect 7026 -1518 7636 -1466
rect 7688 -1468 8248 -1466
rect 7688 -1518 8068 -1468
rect 6466 -1520 8068 -1518
rect 8120 -1470 8248 -1468
rect 8120 -1520 8180 -1470
rect 6466 -1522 8180 -1520
rect 8232 -1522 8248 -1470
rect 6466 -1524 8248 -1522
rect 5799 -1529 8248 -1524
rect 5247 -1541 8248 -1529
rect 5184 -1550 8248 -1541
rect 5194 -1558 5248 -1550
rect 6410 -1560 6470 -1550
rect 6970 -1554 7030 -1550
rect 7102 -1794 7304 -1550
rect 7632 -1554 7692 -1550
rect 8064 -1556 8124 -1550
rect 8176 -1558 8236 -1550
rect 7100 -1806 7304 -1794
rect 4394 -1812 7304 -1806
rect 8868 -1812 8982 -400
rect 9022 -402 9076 -392
rect 9132 -396 9186 -392
rect 4394 -1823 8982 -1812
rect 4394 -1939 7111 -1823
rect 7291 -1868 8982 -1823
rect 7291 -1939 8976 -1868
rect 4394 -1942 8976 -1939
rect 4394 -1968 7302 -1942
rect 4394 -1978 7246 -1968
use sky130_fd_pr__pfet_01v8_GCKZD5  XM1
timestamp 1712816020
transform 1 0 7931 0 1 791
box -479 -419 479 419
use sky130_fd_pr__pfet_01v8_NVWXJJ  XM2
timestamp 1712816020
transform 1 0 4461 0 1 2006
box -385 -544 385 544
use sky130_fd_pr__nfet_01v8_EWGL24  XM3
timestamp 1712816020
transform 1 0 4469 0 1 803
box -375 -525 375 525
use sky130_fd_pr__pfet_01v8_NVWXJJ  XM4
timestamp 1712816020
transform 1 0 5485 0 1 2006
box -385 -544 385 544
use sky130_fd_pr__nfet_01v8_A69A5U  XM5
timestamp 1712816020
transform 1 0 5459 0 1 -159
box -365 -425 365 425
use sky130_fd_pr__pfet_01v8_NVWXJJ  XM6
timestamp 1712816020
transform 1 0 6509 0 1 2008
box -385 -544 385 544
use sky130_fd_pr__pfet_01v8_GCKZD5  XM7
timestamp 1712816020
transform 1 0 5507 0 1 789
box -479 -419 479 419
use sky130_fd_pr__pfet_01v8_GCKZD5  XM8
timestamp 1712816020
transform 1 0 6719 0 1 791
box -479 -419 479 419
use sky130_fd_pr__pfet_01v8_NVWXJJ  XM9
timestamp 1712816020
transform 1 0 7533 0 1 2008
box -385 -544 385 544
use sky130_fd_pr__nfet_01v8_A69A5U  XM10
timestamp 1712816020
transform 1 0 6661 0 1 -161
box -365 -425 365 425
use sky130_fd_pr__nfet_01v8_A69A5U  XM11
timestamp 1712816020
transform 1 0 7879 0 1 -157
box -365 -425 365 425
use sky130_fd_pr__nfet_01v8_EWGL24  XM12
timestamp 1712816020
transform 1 0 5441 0 1 -1225
box -375 -525 375 525
use sky130_fd_pr__nfet_01v8_EWGL24  XM13
timestamp 1712816020
transform 1 0 6657 0 1 -1229
box -375 -525 375 525
use sky130_fd_pr__nfet_01v8_EWGL24  XM14
timestamp 1712816020
transform 1 0 7877 0 1 -1229
box -375 -525 375 525
use sky130_fd_pr__nfet_01v8_ZAY3BZ  XM15
timestamp 1712816020
transform 1 0 8951 0 1 -171
box -253 -425 253 425
use sky130_fd_pr__pfet_01v8_XGJZDL  XM16
timestamp 1712816020
transform 1 0 8977 0 1 803
box -311 -419 311 419
<< labels >>
flabel metal1 s 3508 578 3708 778 0 FreeSans 626 0 0 0 vctrl
port 1 nsew
flabel metal1 s 5948 2734 6148 2934 0 FreeSans 626 0 0 0 VDD
port 2 nsew
flabel metal1 s 7098 -2212 7298 -2012 0 FreeSans 626 0 0 0 VSS
port 3 nsew
flabel metal1 s 9378 234 9578 434 0 FreeSans 626 0 0 0 Osc_out
port 4 nsew
<< end >>
