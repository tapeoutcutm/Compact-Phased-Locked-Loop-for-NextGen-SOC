magic
tech sky130A
magscale 1 2
timestamp 1712816020
<< nwell >>
rect 5986 940 6210 1246
<< pwell >>
rect 6012 604 6162 814
<< psubdiff >>
rect 6038 753 6136 788
rect 6038 719 6069 753
rect 6103 719 6136 753
rect 6038 685 6136 719
rect 6038 651 6069 685
rect 6103 651 6136 685
rect 6038 630 6136 651
<< nsubdiff >>
rect 6036 1156 6138 1198
rect 6036 1122 6067 1156
rect 6101 1122 6138 1156
rect 6036 1088 6138 1122
rect 6036 1054 6067 1088
rect 6101 1054 6138 1088
rect 6036 990 6138 1054
<< psubdiffcont >>
rect 6069 719 6103 753
rect 6069 651 6103 685
<< nsubdiffcont >>
rect 6067 1122 6101 1156
rect 6067 1054 6101 1088
<< locali >>
rect 6036 1166 6138 1198
rect 5672 1156 6138 1166
rect 5944 1128 6067 1156
rect 6036 1122 6067 1128
rect 6101 1122 6138 1156
rect 6036 1088 6138 1122
rect 6036 1054 6067 1088
rect 6101 1054 6138 1088
rect 6036 990 6138 1054
rect 1576 854 1678 920
rect -202 800 -64 834
rect 140 806 178 816
rect 1920 815 1966 832
rect 3370 828 3590 858
rect 140 772 142 806
rect 176 772 178 806
rect 140 762 178 772
rect 1548 804 1586 814
rect 1548 770 1550 804
rect 1584 770 1586 804
rect 1548 760 1586 770
rect 1920 781 1926 815
rect 1960 781 1966 815
rect 1920 764 1966 781
rect 3328 811 3590 828
rect 3328 777 3334 811
rect 3368 802 3590 811
rect 3842 835 3888 852
rect 3368 777 3374 802
rect 3842 801 3848 835
rect 3882 801 3888 835
rect 3842 784 3888 801
rect 5248 831 5294 848
rect 5248 797 5254 831
rect 5288 797 5294 831
rect 5524 816 5702 864
rect 5952 862 6002 886
rect 5834 858 6002 862
rect 5834 824 5960 858
rect 5994 824 6002 858
rect 5834 822 6002 824
rect 5248 780 5294 797
rect 5952 796 6002 822
rect 3328 760 3374 777
rect 6038 753 6136 788
rect 4952 726 4994 730
rect 4952 692 4956 726
rect 4990 692 4994 726
rect 4952 688 4994 692
rect 6038 719 6069 753
rect 6103 719 6136 753
rect 6038 685 6136 719
rect 6038 651 6069 685
rect 6103 651 6136 685
rect 6038 630 6136 651
rect 5918 584 6136 630
<< viali >>
rect -236 800 -202 834
rect 142 772 176 806
rect 1550 770 1584 804
rect 1926 781 1960 815
rect 3334 777 3368 811
rect 3848 801 3882 835
rect 5254 797 5288 831
rect 5392 820 5426 854
rect 5960 824 5994 858
rect 4956 692 4990 726
<< metal1 >>
rect -402 994 -202 1194
rect 0 1096 5948 1192
rect 5948 898 6148 942
rect -397 877 -197 891
rect -397 865 -195 877
rect -397 834 -153 865
rect 3836 852 3894 864
rect 5242 852 5300 860
rect -397 800 -236 834
rect -202 800 -153 834
rect 1914 832 1972 844
rect 3322 832 3380 840
rect -397 771 -153 800
rect 134 816 184 828
rect 1542 816 1592 826
rect 134 806 1592 816
rect 134 772 142 806
rect 176 804 1592 806
rect 176 772 1550 804
rect -397 757 -195 771
rect 134 770 1550 772
rect 1584 770 1592 804
rect 134 760 1592 770
rect -397 691 -197 757
rect 134 750 184 760
rect 1542 748 1592 760
rect 1914 815 3380 832
rect 1914 781 1926 815
rect 1960 811 3380 815
rect 1960 781 3334 811
rect 1914 777 3334 781
rect 3368 777 3380 811
rect 1914 766 3380 777
rect 3836 835 5300 852
rect 3836 801 3848 835
rect 3882 831 5300 835
rect 3882 801 5254 831
rect 3836 797 5254 801
rect 5288 797 5300 831
rect 3836 786 5300 797
rect 3836 772 3894 786
rect 5242 768 5300 786
rect 5380 854 5438 860
rect 5380 820 5392 854
rect 5426 820 5438 854
rect 1914 752 1972 766
rect 3322 748 3380 766
rect 5380 738 5438 820
rect 5946 858 6148 898
rect 5946 824 5960 858
rect 5994 824 6148 858
rect 5946 784 6148 824
rect 5948 742 6148 784
rect 4948 736 5438 738
rect 4940 726 5438 736
rect 4940 692 4956 726
rect 4990 692 5438 726
rect 4940 682 5438 692
rect 4948 680 5438 682
rect 4948 678 5430 680
rect 0 552 6148 648
rect 5948 448 6148 552
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_0
timestamp 1712816020
transform 1 0 -230 0 1 600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_1
timestamp 1712816020
transform 1 0 3434 0 1 600
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1#0  x1
timestamp 1712816020
transform 1 0 -138 0 1 600
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxbp_1#0  x2
timestamp 1712816020
transform 1 0 1644 0 1 600
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxbp_1#0  x3
timestamp 1712816020
transform 1 0 3564 0 1 600
box -38 -48 1786 592
use sky130_fd_sc_hd__inv_2  x4
timestamp 1712816020
transform 1 0 5358 0 1 600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  x5
timestamp 1712816020
transform 1 0 5672 0 1 600
box -38 -48 314 592
<< labels >>
flabel metal1 s -397 691 -197 891 0 FreeSans 626 0 0 0 f0
port 1 nsew
flabel metal1 s -402 994 -202 1194 0 FreeSans 626 0 0 0 VDD
port 2 nsew
flabel metal1 s 5948 742 6148 942 0 FreeSans 626 0 0 0 f0_by_8
port 3 nsew
flabel metal1 s 5948 448 6148 648 0 FreeSans 626 0 0 0 VSS
port 4 nsew
<< end >>
