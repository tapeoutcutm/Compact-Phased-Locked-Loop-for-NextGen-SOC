magic
tech sky130A
magscale 1 2
timestamp 1712816020
<< error_p >>
rect -29 281 29 287
rect -29 247 -17 281
rect -29 241 29 247
rect -125 -247 -67 -241
rect 67 -247 125 -241
rect -125 -281 -113 -247
rect 67 -281 79 -247
rect -125 -287 -67 -281
rect 67 -287 125 -281
<< nwell >>
rect -311 -419 311 419
<< pmos >>
rect -111 -200 -81 200
rect -15 -200 15 200
rect 81 -200 111 200
<< pdiff >>
rect -173 187 -111 200
rect -173 153 -161 187
rect -127 153 -111 187
rect -173 119 -111 153
rect -173 85 -161 119
rect -127 85 -111 119
rect -173 51 -111 85
rect -173 17 -161 51
rect -127 17 -111 51
rect -173 -17 -111 17
rect -173 -51 -161 -17
rect -127 -51 -111 -17
rect -173 -85 -111 -51
rect -173 -119 -161 -85
rect -127 -119 -111 -85
rect -173 -153 -111 -119
rect -173 -187 -161 -153
rect -127 -187 -111 -153
rect -173 -200 -111 -187
rect -81 187 -15 200
rect -81 153 -65 187
rect -31 153 -15 187
rect -81 119 -15 153
rect -81 85 -65 119
rect -31 85 -15 119
rect -81 51 -15 85
rect -81 17 -65 51
rect -31 17 -15 51
rect -81 -17 -15 17
rect -81 -51 -65 -17
rect -31 -51 -15 -17
rect -81 -85 -15 -51
rect -81 -119 -65 -85
rect -31 -119 -15 -85
rect -81 -153 -15 -119
rect -81 -187 -65 -153
rect -31 -187 -15 -153
rect -81 -200 -15 -187
rect 15 187 81 200
rect 15 153 31 187
rect 65 153 81 187
rect 15 119 81 153
rect 15 85 31 119
rect 65 85 81 119
rect 15 51 81 85
rect 15 17 31 51
rect 65 17 81 51
rect 15 -17 81 17
rect 15 -51 31 -17
rect 65 -51 81 -17
rect 15 -85 81 -51
rect 15 -119 31 -85
rect 65 -119 81 -85
rect 15 -153 81 -119
rect 15 -187 31 -153
rect 65 -187 81 -153
rect 15 -200 81 -187
rect 111 187 173 200
rect 111 153 127 187
rect 161 153 173 187
rect 111 119 173 153
rect 111 85 127 119
rect 161 85 173 119
rect 111 51 173 85
rect 111 17 127 51
rect 161 17 173 51
rect 111 -17 173 17
rect 111 -51 127 -17
rect 161 -51 173 -17
rect 111 -85 173 -51
rect 111 -119 127 -85
rect 161 -119 173 -85
rect 111 -153 173 -119
rect 111 -187 127 -153
rect 161 -187 173 -153
rect 111 -200 173 -187
<< pdiffc >>
rect -161 153 -127 187
rect -161 85 -127 119
rect -161 17 -127 51
rect -161 -51 -127 -17
rect -161 -119 -127 -85
rect -161 -187 -127 -153
rect -65 153 -31 187
rect -65 85 -31 119
rect -65 17 -31 51
rect -65 -51 -31 -17
rect -65 -119 -31 -85
rect -65 -187 -31 -153
rect 31 153 65 187
rect 31 85 65 119
rect 31 17 65 51
rect 31 -51 65 -17
rect 31 -119 65 -85
rect 31 -187 65 -153
rect 127 153 161 187
rect 127 85 161 119
rect 127 17 161 51
rect 127 -51 161 -17
rect 127 -119 161 -85
rect 127 -187 161 -153
<< nsubdiff >>
rect -275 349 -153 383
rect -119 349 -85 383
rect -51 349 -17 383
rect 17 349 51 383
rect 85 349 119 383
rect 153 349 275 383
rect -275 255 -241 349
rect 241 255 275 349
rect -275 187 -241 221
rect -275 119 -241 153
rect -275 51 -241 85
rect -275 -17 -241 17
rect -275 -85 -241 -51
rect -275 -153 -241 -119
rect -275 -221 -241 -187
rect 241 187 275 221
rect 241 119 275 153
rect 241 51 275 85
rect 241 -17 275 17
rect 241 -85 275 -51
rect 241 -153 275 -119
rect 241 -221 275 -187
rect -275 -349 -241 -255
rect 241 -349 275 -255
rect -275 -383 -153 -349
rect -119 -383 -85 -349
rect -51 -383 -17 -349
rect 17 -383 51 -349
rect 85 -383 119 -349
rect 153 -383 275 -349
<< nsubdiffcont >>
rect -153 349 -119 383
rect -85 349 -51 383
rect -17 349 17 383
rect 51 349 85 383
rect 119 349 153 383
rect -275 221 -241 255
rect 241 221 275 255
rect -275 153 -241 187
rect -275 85 -241 119
rect -275 17 -241 51
rect -275 -51 -241 -17
rect -275 -119 -241 -85
rect -275 -187 -241 -153
rect 241 153 275 187
rect 241 85 275 119
rect 241 17 275 51
rect 241 -51 275 -17
rect 241 -119 275 -85
rect 241 -187 275 -153
rect -275 -255 -241 -221
rect 241 -255 275 -221
rect -153 -383 -119 -349
rect -85 -383 -51 -349
rect -17 -383 17 -349
rect 51 -383 85 -349
rect 119 -383 153 -349
<< poly >>
rect -33 281 33 297
rect -33 247 -17 281
rect 17 247 33 281
rect -33 231 33 247
rect -111 200 -81 226
rect -15 200 15 231
rect 81 200 111 226
rect -111 -231 -81 -200
rect -15 -226 15 -200
rect 81 -231 111 -200
rect -129 -247 -63 -231
rect -129 -281 -113 -247
rect -79 -281 -63 -247
rect -129 -297 -63 -281
rect 63 -247 129 -231
rect 63 -281 79 -247
rect 113 -281 129 -247
rect 63 -297 129 -281
<< polycont >>
rect -17 247 17 281
rect -113 -281 -79 -247
rect 79 -281 113 -247
<< locali >>
rect -275 349 -153 383
rect -119 349 -85 383
rect -51 349 -17 383
rect 17 349 51 383
rect 85 349 119 383
rect 153 349 275 383
rect -275 255 -241 349
rect -33 247 -17 281
rect 17 247 33 281
rect 241 255 275 349
rect -275 187 -241 221
rect -275 119 -241 153
rect -275 51 -241 85
rect -275 -17 -241 17
rect -275 -85 -241 -51
rect -275 -153 -241 -119
rect -275 -221 -241 -187
rect -161 187 -127 204
rect -161 119 -127 127
rect -161 51 -127 55
rect -161 -55 -127 -51
rect -161 -127 -127 -119
rect -161 -204 -127 -187
rect -65 187 -31 204
rect -65 119 -31 127
rect -65 51 -31 55
rect -65 -55 -31 -51
rect -65 -127 -31 -119
rect -65 -204 -31 -187
rect 31 187 65 204
rect 31 119 65 127
rect 31 51 65 55
rect 31 -55 65 -51
rect 31 -127 65 -119
rect 31 -204 65 -187
rect 127 187 161 204
rect 127 119 161 127
rect 127 51 161 55
rect 127 -55 161 -51
rect 127 -127 161 -119
rect 127 -204 161 -187
rect 241 187 275 221
rect 241 119 275 153
rect 241 51 275 85
rect 241 -17 275 17
rect 241 -85 275 -51
rect 241 -153 275 -119
rect 241 -221 275 -187
rect -275 -349 -241 -255
rect -129 -281 -113 -247
rect -79 -281 -63 -247
rect 63 -281 79 -247
rect 113 -281 129 -247
rect 241 -349 275 -255
rect -275 -383 -153 -349
rect -119 -383 -85 -349
rect -51 -383 -17 -349
rect 17 -383 51 -349
rect 85 -383 119 -349
rect 153 -383 275 -349
<< viali >>
rect -17 247 17 281
rect -161 153 -127 161
rect -161 127 -127 153
rect -161 85 -127 89
rect -161 55 -127 85
rect -161 -17 -127 17
rect -161 -85 -127 -55
rect -161 -89 -127 -85
rect -161 -153 -127 -127
rect -161 -161 -127 -153
rect -65 153 -31 161
rect -65 127 -31 153
rect -65 85 -31 89
rect -65 55 -31 85
rect -65 -17 -31 17
rect -65 -85 -31 -55
rect -65 -89 -31 -85
rect -65 -153 -31 -127
rect -65 -161 -31 -153
rect 31 153 65 161
rect 31 127 65 153
rect 31 85 65 89
rect 31 55 65 85
rect 31 -17 65 17
rect 31 -85 65 -55
rect 31 -89 65 -85
rect 31 -153 65 -127
rect 31 -161 65 -153
rect 127 153 161 161
rect 127 127 161 153
rect 127 85 161 89
rect 127 55 161 85
rect 127 -17 161 17
rect 127 -85 161 -55
rect 127 -89 161 -85
rect 127 -153 161 -127
rect 127 -161 161 -153
rect -113 -281 -79 -247
rect 79 -281 113 -247
<< metal1 >>
rect -29 281 29 287
rect -29 247 -17 281
rect 17 247 29 281
rect -29 241 29 247
rect -167 161 -121 200
rect -167 127 -161 161
rect -127 127 -121 161
rect -167 89 -121 127
rect -167 55 -161 89
rect -127 55 -121 89
rect -167 17 -121 55
rect -167 -17 -161 17
rect -127 -17 -121 17
rect -167 -55 -121 -17
rect -167 -89 -161 -55
rect -127 -89 -121 -55
rect -167 -127 -121 -89
rect -167 -161 -161 -127
rect -127 -161 -121 -127
rect -167 -200 -121 -161
rect -71 161 -25 200
rect -71 127 -65 161
rect -31 127 -25 161
rect -71 89 -25 127
rect -71 55 -65 89
rect -31 55 -25 89
rect -71 17 -25 55
rect -71 -17 -65 17
rect -31 -17 -25 17
rect -71 -55 -25 -17
rect -71 -89 -65 -55
rect -31 -89 -25 -55
rect -71 -127 -25 -89
rect -71 -161 -65 -127
rect -31 -161 -25 -127
rect -71 -200 -25 -161
rect 25 161 71 200
rect 25 127 31 161
rect 65 127 71 161
rect 25 89 71 127
rect 25 55 31 89
rect 65 55 71 89
rect 25 17 71 55
rect 25 -17 31 17
rect 65 -17 71 17
rect 25 -55 71 -17
rect 25 -89 31 -55
rect 65 -89 71 -55
rect 25 -127 71 -89
rect 25 -161 31 -127
rect 65 -161 71 -127
rect 25 -200 71 -161
rect 121 161 167 200
rect 121 127 127 161
rect 161 127 167 161
rect 121 89 167 127
rect 121 55 127 89
rect 161 55 167 89
rect 121 17 167 55
rect 121 -17 127 17
rect 161 -17 167 17
rect 121 -55 167 -17
rect 121 -89 127 -55
rect 161 -89 167 -55
rect 121 -127 167 -89
rect 121 -161 127 -127
rect 161 -161 167 -127
rect 121 -200 167 -161
rect -125 -247 -67 -241
rect -125 -281 -113 -247
rect -79 -281 -67 -247
rect -125 -287 -67 -281
rect 67 -247 125 -241
rect 67 -281 79 -247
rect 113 -281 125 -247
rect 67 -287 125 -281
<< properties >>
string FIXED_BBOX -258 -366 258 366
<< end >>
