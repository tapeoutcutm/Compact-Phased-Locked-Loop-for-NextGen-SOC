magic
tech sky130A
magscale 1 2
timestamp 1712816020
<< error_p >>
rect 19 297 77 303
rect 19 263 31 297
rect 19 257 77 263
rect -77 -263 -19 -257
rect -77 -297 -65 -263
rect -77 -303 -19 -297
<< pwell >>
rect -253 -425 253 425
<< nmos >>
rect -63 -225 -33 225
rect 33 -225 63 225
<< ndiff >>
rect -125 187 -63 225
rect -125 153 -113 187
rect -79 153 -63 187
rect -125 119 -63 153
rect -125 85 -113 119
rect -79 85 -63 119
rect -125 51 -63 85
rect -125 17 -113 51
rect -79 17 -63 51
rect -125 -17 -63 17
rect -125 -51 -113 -17
rect -79 -51 -63 -17
rect -125 -85 -63 -51
rect -125 -119 -113 -85
rect -79 -119 -63 -85
rect -125 -153 -63 -119
rect -125 -187 -113 -153
rect -79 -187 -63 -153
rect -125 -225 -63 -187
rect -33 187 33 225
rect -33 153 -17 187
rect 17 153 33 187
rect -33 119 33 153
rect -33 85 -17 119
rect 17 85 33 119
rect -33 51 33 85
rect -33 17 -17 51
rect 17 17 33 51
rect -33 -17 33 17
rect -33 -51 -17 -17
rect 17 -51 33 -17
rect -33 -85 33 -51
rect -33 -119 -17 -85
rect 17 -119 33 -85
rect -33 -153 33 -119
rect -33 -187 -17 -153
rect 17 -187 33 -153
rect -33 -225 33 -187
rect 63 187 125 225
rect 63 153 79 187
rect 113 153 125 187
rect 63 119 125 153
rect 63 85 79 119
rect 113 85 125 119
rect 63 51 125 85
rect 63 17 79 51
rect 113 17 125 51
rect 63 -17 125 17
rect 63 -51 79 -17
rect 113 -51 125 -17
rect 63 -85 125 -51
rect 63 -119 79 -85
rect 113 -119 125 -85
rect 63 -153 125 -119
rect 63 -187 79 -153
rect 113 -187 125 -153
rect 63 -225 125 -187
<< ndiffc >>
rect -113 153 -79 187
rect -113 85 -79 119
rect -113 17 -79 51
rect -113 -51 -79 -17
rect -113 -119 -79 -85
rect -113 -187 -79 -153
rect -17 153 17 187
rect -17 85 17 119
rect -17 17 17 51
rect -17 -51 17 -17
rect -17 -119 17 -85
rect -17 -187 17 -153
rect 79 153 113 187
rect 79 85 113 119
rect 79 17 113 51
rect 79 -51 113 -17
rect 79 -119 113 -85
rect 79 -187 113 -153
<< psubdiff >>
rect -227 365 -119 399
rect -85 365 -51 399
rect -17 365 17 399
rect 51 365 85 399
rect 119 365 227 399
rect -227 289 -193 365
rect -227 221 -193 255
rect 193 289 227 365
rect -227 153 -193 187
rect -227 85 -193 119
rect -227 17 -193 51
rect -227 -51 -193 -17
rect -227 -119 -193 -85
rect -227 -187 -193 -153
rect -227 -255 -193 -221
rect 193 221 227 255
rect 193 153 227 187
rect 193 85 227 119
rect 193 17 227 51
rect 193 -51 227 -17
rect 193 -119 227 -85
rect 193 -187 227 -153
rect -227 -365 -193 -289
rect 193 -255 227 -221
rect 193 -365 227 -289
rect -227 -399 -119 -365
rect -85 -399 -51 -365
rect -17 -399 17 -365
rect 51 -399 85 -365
rect 119 -399 227 -365
<< psubdiffcont >>
rect -119 365 -85 399
rect -51 365 -17 399
rect 17 365 51 399
rect 85 365 119 399
rect -227 255 -193 289
rect 193 255 227 289
rect -227 187 -193 221
rect -227 119 -193 153
rect -227 51 -193 85
rect -227 -17 -193 17
rect -227 -85 -193 -51
rect -227 -153 -193 -119
rect -227 -221 -193 -187
rect 193 187 227 221
rect 193 119 227 153
rect 193 51 227 85
rect 193 -17 227 17
rect 193 -85 227 -51
rect 193 -153 227 -119
rect 193 -221 227 -187
rect -227 -289 -193 -255
rect 193 -289 227 -255
rect -119 -399 -85 -365
rect -51 -399 -17 -365
rect 17 -399 51 -365
rect 85 -399 119 -365
<< poly >>
rect 15 297 81 313
rect 15 263 31 297
rect 65 263 81 297
rect -63 225 -33 251
rect 15 247 81 263
rect 33 225 63 247
rect -63 -247 -33 -225
rect -81 -263 -15 -247
rect 33 -251 63 -225
rect -81 -297 -65 -263
rect -31 -297 -15 -263
rect -81 -313 -15 -297
<< polycont >>
rect 31 263 65 297
rect -65 -297 -31 -263
<< locali >>
rect -227 365 -119 399
rect -85 365 -51 399
rect -17 365 17 399
rect 51 365 85 399
rect 119 365 227 399
rect -227 289 -193 365
rect 15 263 31 297
rect 65 263 81 297
rect 193 289 227 365
rect -227 221 -193 255
rect -227 153 -193 187
rect -227 85 -193 119
rect -227 17 -193 51
rect -227 -51 -193 -17
rect -227 -119 -193 -85
rect -227 -187 -193 -153
rect -227 -255 -193 -221
rect -113 197 -79 229
rect -113 125 -79 153
rect -113 53 -79 85
rect -113 -17 -79 17
rect -113 -85 -79 -53
rect -113 -153 -79 -125
rect -113 -229 -79 -197
rect -17 197 17 229
rect -17 125 17 153
rect -17 53 17 85
rect -17 -17 17 17
rect -17 -85 17 -53
rect -17 -153 17 -125
rect -17 -229 17 -197
rect 79 197 113 229
rect 79 125 113 153
rect 79 53 113 85
rect 79 -17 113 17
rect 79 -85 113 -53
rect 79 -153 113 -125
rect 79 -229 113 -197
rect 193 221 227 255
rect 193 153 227 187
rect 193 85 227 119
rect 193 17 227 51
rect 193 -51 227 -17
rect 193 -119 227 -85
rect 193 -187 227 -153
rect 193 -255 227 -221
rect -227 -365 -193 -289
rect -81 -297 -65 -263
rect -31 -297 -15 -263
rect 193 -365 227 -289
rect -227 -399 -119 -365
rect -85 -399 -51 -365
rect -17 -399 17 -365
rect 51 -399 85 -365
rect 119 -399 227 -365
<< viali >>
rect 31 263 65 297
rect -113 187 -79 197
rect -113 163 -79 187
rect -113 119 -79 125
rect -113 91 -79 119
rect -113 51 -79 53
rect -113 19 -79 51
rect -113 -51 -79 -19
rect -113 -53 -79 -51
rect -113 -119 -79 -91
rect -113 -125 -79 -119
rect -113 -187 -79 -163
rect -113 -197 -79 -187
rect -17 187 17 197
rect -17 163 17 187
rect -17 119 17 125
rect -17 91 17 119
rect -17 51 17 53
rect -17 19 17 51
rect -17 -51 17 -19
rect -17 -53 17 -51
rect -17 -119 17 -91
rect -17 -125 17 -119
rect -17 -187 17 -163
rect -17 -197 17 -187
rect 79 187 113 197
rect 79 163 113 187
rect 79 119 113 125
rect 79 91 113 119
rect 79 51 113 53
rect 79 19 113 51
rect 79 -51 113 -19
rect 79 -53 113 -51
rect 79 -119 113 -91
rect 79 -125 113 -119
rect 79 -187 113 -163
rect 79 -197 113 -187
rect -65 -297 -31 -263
<< metal1 >>
rect 19 297 77 303
rect 19 263 31 297
rect 65 263 77 297
rect 19 257 77 263
rect -119 197 -73 225
rect -119 163 -113 197
rect -79 163 -73 197
rect -119 125 -73 163
rect -119 91 -113 125
rect -79 91 -73 125
rect -119 53 -73 91
rect -119 19 -113 53
rect -79 19 -73 53
rect -119 -19 -73 19
rect -119 -53 -113 -19
rect -79 -53 -73 -19
rect -119 -91 -73 -53
rect -119 -125 -113 -91
rect -79 -125 -73 -91
rect -119 -163 -73 -125
rect -119 -197 -113 -163
rect -79 -197 -73 -163
rect -119 -225 -73 -197
rect -23 197 23 225
rect -23 163 -17 197
rect 17 163 23 197
rect -23 125 23 163
rect -23 91 -17 125
rect 17 91 23 125
rect -23 53 23 91
rect -23 19 -17 53
rect 17 19 23 53
rect -23 -19 23 19
rect -23 -53 -17 -19
rect 17 -53 23 -19
rect -23 -91 23 -53
rect -23 -125 -17 -91
rect 17 -125 23 -91
rect -23 -163 23 -125
rect -23 -197 -17 -163
rect 17 -197 23 -163
rect -23 -225 23 -197
rect 73 197 119 225
rect 73 163 79 197
rect 113 163 119 197
rect 73 125 119 163
rect 73 91 79 125
rect 113 91 119 125
rect 73 53 119 91
rect 73 19 79 53
rect 113 19 119 53
rect 73 -19 119 19
rect 73 -53 79 -19
rect 113 -53 119 -19
rect 73 -91 119 -53
rect 73 -125 79 -91
rect 113 -125 119 -91
rect 73 -163 119 -125
rect 73 -197 79 -163
rect 113 -197 119 -163
rect 73 -225 119 -197
rect -77 -263 -19 -257
rect -77 -297 -65 -263
rect -31 -297 -19 -263
rect -77 -303 -19 -297
<< properties >>
string FIXED_BBOX -210 -382 210 382
<< end >>
