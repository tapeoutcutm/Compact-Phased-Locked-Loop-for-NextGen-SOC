magic
tech sky130A
magscale 1 2
timestamp 1712816020
<< nwell >>
rect -396 -319 396 319
<< pmos >>
rect -200 -100 200 100
<< pdiff >>
rect -258 85 -200 100
rect -258 51 -246 85
rect -212 51 -200 85
rect -258 17 -200 51
rect -258 -17 -246 17
rect -212 -17 -200 17
rect -258 -51 -200 -17
rect -258 -85 -246 -51
rect -212 -85 -200 -51
rect -258 -100 -200 -85
rect 200 85 258 100
rect 200 51 212 85
rect 246 51 258 85
rect 200 17 258 51
rect 200 -17 212 17
rect 246 -17 258 17
rect 200 -51 258 -17
rect 200 -85 212 -51
rect 246 -85 258 -51
rect 200 -100 258 -85
<< pdiffc >>
rect -246 51 -212 85
rect -246 -17 -212 17
rect -246 -85 -212 -51
rect 212 51 246 85
rect 212 -17 246 17
rect 212 -85 246 -51
<< nsubdiff >>
rect -360 249 -255 283
rect -221 249 -187 283
rect -153 249 -119 283
rect -85 249 -51 283
rect -17 249 17 283
rect 51 249 85 283
rect 119 249 153 283
rect 187 249 221 283
rect 255 249 360 283
rect -360 187 -326 249
rect -360 119 -326 153
rect 326 187 360 249
rect 326 119 360 153
rect -360 51 -326 85
rect -360 -17 -326 17
rect -360 -85 -326 -51
rect 326 51 360 85
rect 326 -17 360 17
rect 326 -85 360 -51
rect -360 -153 -326 -119
rect -360 -249 -326 -187
rect 326 -153 360 -119
rect 326 -249 360 -187
rect -360 -283 -255 -249
rect -221 -283 -187 -249
rect -153 -283 -119 -249
rect -85 -283 -51 -249
rect -17 -283 17 -249
rect 51 -283 85 -249
rect 119 -283 153 -249
rect 187 -283 221 -249
rect 255 -283 360 -249
<< nsubdiffcont >>
rect -255 249 -221 283
rect -187 249 -153 283
rect -119 249 -85 283
rect -51 249 -17 283
rect 17 249 51 283
rect 85 249 119 283
rect 153 249 187 283
rect 221 249 255 283
rect -360 153 -326 187
rect -360 85 -326 119
rect 326 153 360 187
rect -360 17 -326 51
rect -360 -51 -326 -17
rect -360 -119 -326 -85
rect 326 85 360 119
rect 326 17 360 51
rect 326 -51 360 -17
rect -360 -187 -326 -153
rect 326 -119 360 -85
rect 326 -187 360 -153
rect -255 -283 -221 -249
rect -187 -283 -153 -249
rect -119 -283 -85 -249
rect -51 -283 -17 -249
rect 17 -283 51 -249
rect 85 -283 119 -249
rect 153 -283 187 -249
rect 221 -283 255 -249
<< poly >>
rect -200 181 200 197
rect -200 147 -153 181
rect -119 147 -85 181
rect -51 147 -17 181
rect 17 147 51 181
rect 85 147 119 181
rect 153 147 200 181
rect -200 100 200 147
rect -200 -147 200 -100
rect -200 -181 -153 -147
rect -119 -181 -85 -147
rect -51 -181 -17 -147
rect 17 -181 51 -147
rect 85 -181 119 -147
rect 153 -181 200 -147
rect -200 -197 200 -181
<< polycont >>
rect -153 147 -119 181
rect -85 147 -51 181
rect -17 147 17 181
rect 51 147 85 181
rect 119 147 153 181
rect -153 -181 -119 -147
rect -85 -181 -51 -147
rect -17 -181 17 -147
rect 51 -181 85 -147
rect 119 -181 153 -147
<< locali >>
rect -360 249 -255 283
rect -221 249 -187 283
rect -153 249 -119 283
rect -85 249 -51 283
rect -17 249 17 283
rect 51 249 85 283
rect 119 249 153 283
rect 187 249 221 283
rect 255 249 360 283
rect -360 187 -326 249
rect 326 187 360 249
rect -360 119 -326 153
rect -200 147 -161 181
rect -119 147 -89 181
rect -51 147 -17 181
rect 17 147 51 181
rect 89 147 119 181
rect 161 147 200 181
rect 326 119 360 153
rect -360 51 -326 85
rect -360 -17 -326 17
rect -360 -85 -326 -51
rect -246 85 -212 104
rect -246 17 -212 19
rect -246 -19 -212 -17
rect -246 -104 -212 -85
rect 212 85 246 104
rect 212 17 246 19
rect 212 -19 246 -17
rect 212 -104 246 -85
rect 326 51 360 85
rect 326 -17 360 17
rect 326 -85 360 -51
rect -360 -153 -326 -119
rect -200 -181 -161 -147
rect -119 -181 -89 -147
rect -51 -181 -17 -147
rect 17 -181 51 -147
rect 89 -181 119 -147
rect 161 -181 200 -147
rect 326 -153 360 -119
rect -360 -249 -326 -187
rect 326 -249 360 -187
rect -360 -283 -255 -249
rect -221 -283 -187 -249
rect -153 -283 -119 -249
rect -85 -283 -51 -249
rect -17 -283 17 -249
rect 51 -283 85 -249
rect 119 -283 153 -249
rect 187 -283 221 -249
rect 255 -283 360 -249
<< viali >>
rect -161 147 -153 181
rect -153 147 -127 181
rect -89 147 -85 181
rect -85 147 -55 181
rect -17 147 17 181
rect 55 147 85 181
rect 85 147 89 181
rect 127 147 153 181
rect 153 147 161 181
rect -246 51 -212 53
rect -246 19 -212 51
rect -246 -51 -212 -19
rect -246 -53 -212 -51
rect 212 51 246 53
rect 212 19 246 51
rect 212 -51 246 -19
rect 212 -53 246 -51
rect -161 -181 -153 -147
rect -153 -181 -127 -147
rect -89 -181 -85 -147
rect -85 -181 -55 -147
rect -17 -181 17 -147
rect 55 -181 85 -147
rect 85 -181 89 -147
rect 127 -181 153 -147
rect 153 -181 161 -147
<< metal1 >>
rect -196 181 196 187
rect -196 147 -161 181
rect -127 147 -89 181
rect -55 147 -17 181
rect 17 147 55 181
rect 89 147 127 181
rect 161 147 196 181
rect -196 141 196 147
rect -252 53 -206 100
rect -252 19 -246 53
rect -212 19 -206 53
rect -252 -19 -206 19
rect -252 -53 -246 -19
rect -212 -53 -206 -19
rect -252 -100 -206 -53
rect 206 53 252 100
rect 206 19 212 53
rect 246 19 252 53
rect 206 -19 252 19
rect 206 -53 212 -19
rect 246 -53 252 -19
rect 206 -100 252 -53
rect -196 -147 196 -141
rect -196 -181 -161 -147
rect -127 -181 -89 -147
rect -55 -181 -17 -147
rect 17 -181 55 -147
rect 89 -181 127 -147
rect 161 -181 196 -147
rect -196 -187 196 -181
<< properties >>
string FIXED_BBOX -343 -266 343 266
<< end >>
