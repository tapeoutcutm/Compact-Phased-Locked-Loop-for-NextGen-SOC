magic
tech sky130A
magscale 1 2
timestamp 1712557532
<< metal1 >>
rect 8414 44658 8424 44862
rect 8724 44658 8734 44862
rect 9086 44672 9096 44736
rect 9668 44672 9678 44736
rect 1540 44426 1772 44430
rect 1348 44262 1358 44426
rect 1962 44262 1972 44426
rect 1540 42396 1772 44262
rect 6180 42866 6190 43086
rect 6324 42866 6334 43086
rect 8622 42878 8682 44658
rect 9096 43298 9156 44672
rect 10384 44242 12680 44272
rect 10384 44212 12168 44242
rect 8868 43190 8878 43298
rect 9158 43190 9168 43298
rect 9372 42950 9382 43524
rect 9476 42950 9486 43524
rect 8814 42544 8824 42832
rect 9282 42544 9292 42832
rect 1828 41812 2398 42284
rect 1814 41312 1824 41812
rect 2442 41312 2452 41812
rect 4392 41758 4592 41764
rect 3844 41376 3854 41758
rect 5060 41376 5070 41758
rect 4392 40624 4592 41376
rect 9392 41158 9452 42950
rect 6192 41098 9452 41158
rect 6192 40676 6252 41098
rect 10444 40766 10552 44212
rect 12148 44208 12168 44212
rect 12150 44178 12168 44208
rect 12650 44208 12680 44242
rect 12650 44178 12660 44208
rect 10992 43728 11002 44052
rect 11228 43728 11238 44052
rect 15906 43784 21964 43892
rect 22240 43784 22250 43892
rect 27996 43844 28006 44402
rect 28126 43844 28136 44402
rect 15524 42752 15534 43530
rect 15676 42752 15686 43530
rect 25676 43412 25860 43426
rect 25676 43260 25692 43412
rect 25844 43260 26502 43412
rect 25676 43246 25860 43260
rect 21276 42700 21614 42762
rect 10832 42368 10842 42578
rect 11122 42368 11132 42578
rect 15396 42472 15402 42640
rect 15570 42622 15576 42640
rect 21276 42622 21316 42700
rect 15570 42490 21316 42622
rect 15570 42472 15576 42490
rect 21276 42474 21316 42490
rect 21534 42474 21614 42700
rect 21276 42448 21614 42474
rect 8620 40658 10552 40766
rect 1600 39960 1610 40558
rect 1772 40260 1782 40558
rect 11280 40412 11480 42238
rect 16424 41332 16434 41800
rect 16798 41332 16808 41800
rect 1772 40060 2154 40260
rect 1772 39960 1808 40060
rect 1608 39956 1808 39960
rect 11106 39912 11116 40412
rect 11616 39912 11626 40412
rect 4386 39792 10088 39806
rect 4386 39606 9820 39792
rect 9810 39320 9820 39606
rect 10060 39606 10088 39792
rect 16492 39640 16692 41332
rect 16912 40746 16922 41242
rect 17046 40942 17056 41242
rect 22998 41134 23008 41828
rect 23462 41134 23472 41828
rect 17086 40942 17274 40986
rect 17046 40786 17274 40942
rect 17046 40746 17086 40786
rect 23400 40784 23410 40998
rect 23676 40784 23686 40998
rect 16918 40742 17086 40746
rect 17118 40416 17318 40686
rect 25954 40576 25964 40982
rect 26184 40722 26194 40982
rect 26184 40578 26494 40722
rect 26184 40576 26194 40578
rect 17072 39908 17082 40416
rect 17434 39908 17444 40416
rect 10060 39320 10070 39606
rect 16492 39440 21882 39640
rect 18856 38902 18866 39102
rect 19066 38902 19076 39102
rect 22142 38884 22152 39108
rect 22326 38884 22336 39108
rect 18674 37126 18684 37326
rect 18884 37126 18924 37326
rect 22128 37160 22138 37362
rect 22322 37160 22332 37362
rect 9768 36676 9778 37028
rect 10138 36954 10148 37028
rect 10138 36752 19303 36954
rect 10138 36676 10148 36752
rect 27230 36622 27240 37382
rect 27578 36622 27588 37382
rect 9760 35400 9770 36320
rect 10488 36136 10498 36320
rect 25014 36282 25024 36500
rect 25892 36486 25902 36500
rect 25892 36286 26528 36486
rect 28028 36408 28096 43844
rect 26876 36340 28096 36408
rect 25892 36282 25902 36286
rect 10488 36128 26530 36136
rect 10488 36120 27602 36128
rect 10488 36010 27608 36120
rect 10488 35536 26530 36010
rect 27598 35632 27608 36010
rect 10488 35400 10498 35536
rect 22610 6340 22620 6630
rect 23638 6340 23648 6630
rect 23006 5926 23284 6340
rect 27358 4602 27368 4896
rect 27642 4602 27652 4896
rect 25364 3702 25374 4048
rect 25686 3702 25696 4048
rect 19316 3412 19326 3630
rect 19776 3412 19786 3630
rect 29440 3316 29746 3350
rect 29440 3084 29452 3316
rect 29660 3084 29746 3316
rect 29440 3070 29746 3084
rect 31124 3288 31182 3300
rect 31124 3022 31166 3288
rect 31408 3022 31418 3288
rect 31124 3008 31182 3022
rect 29386 2184 29396 2456
rect 29608 2184 29618 2456
rect 21858 694 22086 1184
rect 21680 526 21690 694
rect 22182 526 22192 694
<< via1 >>
rect 8424 44658 8724 44862
rect 9096 44672 9668 44736
rect 1358 44262 1962 44426
rect 6190 42866 6324 43086
rect 8878 43190 9158 43298
rect 9382 42950 9476 43524
rect 8824 42544 9282 42832
rect 1824 41312 2442 41812
rect 3854 41376 5060 41758
rect 12168 44178 12650 44242
rect 11002 43728 11228 44052
rect 21964 43784 22240 43892
rect 28006 43844 28126 44402
rect 15534 42752 15676 43530
rect 25692 43260 25844 43412
rect 10842 42368 11122 42578
rect 15402 42472 15570 42640
rect 21316 42474 21534 42700
rect 1610 39960 1772 40558
rect 16434 41332 16798 41800
rect 11116 39912 11616 40412
rect 9820 39320 10060 39792
rect 16922 40746 17046 41242
rect 23008 41134 23462 41828
rect 23410 40784 23676 40998
rect 25964 40576 26184 40982
rect 17082 39908 17434 40416
rect 18866 38902 19066 39102
rect 22152 38884 22326 39108
rect 18684 37126 18884 37326
rect 22138 37160 22322 37362
rect 9778 36676 10138 37028
rect 27240 36622 27578 37382
rect 9770 35400 10488 36320
rect 25024 36282 25892 36500
rect 26530 35632 27598 36010
rect 22620 6340 23638 6630
rect 27368 4602 27642 4896
rect 25374 3702 25686 4048
rect 19326 3412 19776 3630
rect 29452 3084 29660 3316
rect 31166 3022 31408 3288
rect 29396 2184 29608 2456
rect 21690 526 22182 694
<< metal2 >>
rect 8424 44862 8724 44872
rect 9096 44736 9668 44746
rect 9096 44662 9668 44672
rect 8424 44648 8724 44658
rect 9304 44594 10148 44604
rect 9304 44514 10148 44524
rect 1358 44426 1962 44436
rect 1358 44252 1962 44262
rect 9394 43534 9454 44514
rect 28006 44402 28126 44412
rect 12168 44242 12650 44252
rect 12168 44168 12650 44178
rect 11002 44052 11228 44062
rect 21964 43892 22240 43902
rect 28006 43834 28126 43844
rect 21964 43774 22240 43784
rect 11002 43718 11228 43728
rect 9382 43524 9476 43534
rect 8878 43298 9158 43308
rect 8878 43180 9158 43190
rect 6190 43086 6324 43096
rect 9382 42940 9476 42950
rect 15534 43530 15676 43540
rect 6190 42856 6324 42866
rect 9782 42874 10122 42884
rect 8824 42832 9282 42842
rect 9282 42544 9782 42824
rect 8824 42542 9782 42544
rect 8824 42534 9282 42542
rect 25692 43412 25844 43422
rect 25692 43250 25844 43260
rect 15534 42742 15676 42752
rect 21300 42700 21558 42732
rect 15402 42640 15570 42646
rect 9782 42428 10122 42438
rect 10842 42578 11122 42588
rect 15402 42466 15570 42472
rect 21300 42474 21316 42700
rect 21534 42474 21558 42700
rect 21300 42454 21558 42474
rect 10842 42358 11122 42368
rect 16282 42000 17136 42010
rect 1622 41922 16282 41982
rect 1622 40568 1682 41922
rect 16282 41904 17136 41914
rect 23008 41828 23462 41838
rect 1824 41812 2442 41822
rect 16434 41800 16798 41810
rect 3854 41758 5060 41768
rect 3854 41366 5060 41376
rect 16434 41322 16798 41332
rect 1824 41302 2442 41312
rect 16922 41242 17046 41252
rect 23008 41124 23462 41134
rect 23410 40998 23676 41008
rect 23410 40774 23676 40784
rect 25964 40982 26184 40992
rect 16922 40736 17046 40746
rect 1610 40558 1772 40568
rect 25964 40566 26184 40576
rect 1610 39950 1772 39960
rect 11116 40412 11616 40422
rect 11116 39902 11616 39912
rect 17082 40416 17434 40426
rect 17082 39898 17434 39908
rect 9820 39792 10060 39802
rect 9820 39310 10060 39320
rect 18866 39102 19066 39112
rect 18866 38892 19066 38902
rect 22152 39108 22326 39118
rect 22152 38874 22326 38884
rect 27240 37382 27578 37392
rect 22138 37362 22322 37372
rect 18684 37326 18884 37336
rect 22138 37150 22322 37160
rect 18684 37116 18884 37126
rect 9778 37028 10138 37038
rect 9778 36666 10138 36676
rect 27240 36612 27578 36622
rect 25024 36500 25892 36510
rect 9770 36320 10488 36330
rect 25024 36272 25892 36282
rect 26530 36120 27598 36130
rect 26530 35622 27598 35632
rect 9770 35390 10488 35400
rect 202 6768 1016 6778
rect 22620 6630 23638 6640
rect 1016 6345 22620 6599
rect 23638 6596 28415 6599
rect 23638 6345 28426 6596
rect 22620 6330 23638 6340
rect 202 6072 1016 6082
rect 28036 5612 28426 6345
rect 27368 4896 27642 4906
rect 27368 4592 27642 4602
rect 25374 4048 25686 4058
rect 25374 3692 25686 3702
rect 19326 3630 19776 3640
rect 19326 3402 19776 3412
rect 29452 3316 29660 3326
rect 29452 3074 29660 3084
rect 31166 3288 31408 3298
rect 31166 3012 31408 3022
rect 9794 1482 10588 1492
rect 9794 1026 10588 1036
rect 10332 678 10484 1026
rect 21690 694 22182 704
rect 10332 526 21690 678
rect 27588 678 27740 2776
rect 29396 2456 29608 2466
rect 29396 2174 29608 2184
rect 22182 526 27744 678
rect 21690 516 22182 526
<< via2 >>
rect 8424 44658 8724 44862
rect 9096 44672 9668 44736
rect 9304 44524 10148 44594
rect 1358 44262 1962 44426
rect 12168 44178 12650 44242
rect 11002 43728 11228 44052
rect 21964 43784 22240 43892
rect 28006 43844 28126 44402
rect 8878 43190 9158 43298
rect 6190 42866 6324 43086
rect 9782 42438 10122 42874
rect 15534 42752 15676 43530
rect 25692 43260 25844 43412
rect 10842 42368 11122 42578
rect 21316 42474 21534 42700
rect 16282 41914 17136 42000
rect 1824 41312 2442 41812
rect 3854 41376 5060 41758
rect 16434 41332 16798 41800
rect 16922 40746 17046 41242
rect 23008 41134 23462 41828
rect 23410 40784 23676 40998
rect 25964 40576 26184 40982
rect 11116 39912 11616 40412
rect 17082 39908 17434 40416
rect 9820 39320 10060 39792
rect 18866 38902 19066 39102
rect 22152 38884 22326 39108
rect 18684 37126 18884 37326
rect 22138 37160 22322 37362
rect 9778 36676 10138 37028
rect 27240 36622 27578 37382
rect 9770 35400 10488 36320
rect 25024 36282 25892 36500
rect 26530 36010 27598 36120
rect 26530 35632 27598 36010
rect 202 6082 1016 6768
rect 27368 4602 27642 4896
rect 25374 3702 25686 4048
rect 19326 3412 19776 3630
rect 29452 3084 29660 3316
rect 31166 3022 31408 3288
rect 9794 1036 10588 1482
rect 29396 2184 29608 2456
<< metal3 >>
rect 13636 44874 13646 44924
rect 8412 44862 13646 44874
rect 8412 44814 8424 44862
rect 8414 44658 8424 44814
rect 8724 44824 13646 44862
rect 14104 44824 14114 44924
rect 16620 44858 16684 44864
rect 8724 44814 14110 44824
rect 8724 44658 8734 44814
rect 16684 44796 25902 44856
rect 16620 44788 16684 44794
rect 14322 44760 14858 44784
rect 14322 44752 14342 44760
rect 9076 44736 14342 44752
rect 9076 44692 9096 44736
rect 9086 44672 9096 44692
rect 9668 44692 14342 44736
rect 14844 44692 14858 44760
rect 15874 44692 15938 44698
rect 9668 44672 9678 44692
rect 9086 44667 9678 44672
rect 8414 44653 8734 44658
rect 10148 44612 13036 44632
rect 10092 44599 13036 44612
rect 9294 44594 13036 44599
rect 790 44518 796 44582
rect 860 44518 866 44582
rect 9294 44524 9304 44594
rect 10148 44572 13036 44594
rect 10148 44524 10290 44572
rect 13026 44568 13036 44572
rect 13474 44568 13484 44632
rect 25628 44690 25638 44692
rect 15938 44630 25638 44690
rect 15874 44622 15938 44628
rect 9294 44519 10290 44524
rect 798 43702 858 44518
rect 10092 44512 10290 44519
rect 12194 44506 12258 44510
rect 12184 44504 12258 44506
rect 12184 44500 12194 44504
rect 12860 44502 12866 44504
rect 12258 44442 12866 44502
rect 12860 44440 12866 44442
rect 12930 44440 12936 44504
rect 25628 44478 25638 44630
rect 25752 44478 25762 44692
rect 25892 44666 25902 44796
rect 26022 44666 26032 44856
rect 12248 44436 12258 44440
rect 12184 44434 12258 44436
rect 1348 44426 1972 44431
rect 12184 44430 12248 44434
rect 1348 44412 1358 44426
rect 1332 44352 1358 44412
rect 1348 44262 1358 44352
rect 1962 44370 1972 44426
rect 27222 44414 27378 44426
rect 27222 44370 27292 44414
rect 1962 44350 27292 44370
rect 27356 44350 27378 44414
rect 1962 44310 27378 44350
rect 1962 44262 1972 44310
rect 27222 44306 27378 44310
rect 27996 44402 28136 44407
rect 1348 44257 1972 44262
rect 3360 44096 3424 44102
rect 5200 44094 5210 44244
rect 3424 44034 5210 44094
rect 3360 44026 3424 44032
rect 5200 44020 5210 44034
rect 5282 44020 5292 44244
rect 12158 44242 12660 44247
rect 12158 44178 12168 44242
rect 12650 44178 12660 44242
rect 12158 44173 12660 44178
rect 10992 44052 11238 44057
rect 4470 43764 4476 43828
rect 4540 43826 4546 43828
rect 9792 43826 9802 43864
rect 4540 43766 9802 43826
rect 4540 43764 4546 43766
rect 9792 43702 9802 43766
rect 798 43642 9802 43702
rect 9792 43624 9802 43642
rect 10098 43624 10108 43864
rect 10992 43728 11002 44052
rect 11228 43728 11238 44052
rect 21954 43892 22250 43897
rect 21954 43784 21964 43892
rect 22240 43784 22250 43892
rect 27996 43844 28006 44402
rect 28126 43844 28136 44402
rect 27996 43839 28136 43844
rect 21954 43779 22250 43784
rect 10992 43723 11238 43728
rect 15524 43530 15686 43535
rect 8868 43298 9168 43303
rect 8868 43250 8878 43298
rect 6226 43190 8878 43250
rect 9158 43190 9168 43298
rect 6226 43091 6286 43190
rect 8868 43185 9168 43190
rect 6180 43086 6334 43091
rect 6180 42866 6190 43086
rect 6324 42866 6334 43086
rect 6180 42861 6334 42866
rect 9772 42874 10132 42879
rect 9772 42438 9782 42874
rect 10122 42438 10132 42874
rect 15524 42752 15534 43530
rect 15676 42752 15686 43530
rect 25682 43412 25854 43417
rect 25682 43260 25692 43412
rect 25844 43260 25854 43412
rect 25682 43255 25854 43260
rect 15524 42747 15686 42752
rect 9772 42433 10132 42438
rect 10832 42578 11132 42583
rect 10832 42368 10842 42578
rect 11122 42368 11132 42578
rect 10832 42363 11132 42368
rect 8533 41822 9031 41827
rect 15542 41824 15674 42747
rect 21306 42700 21544 42705
rect 21306 42474 21316 42700
rect 21534 42474 21544 42700
rect 21306 42469 21544 42474
rect 24200 42428 24376 42442
rect 23910 42384 24076 42398
rect 19166 42374 19316 42384
rect 15764 42337 15904 42352
rect 17712 42341 17808 42352
rect 17712 42337 17725 42341
rect 15764 42335 17725 42337
rect 15764 42271 15776 42335
rect 15840 42277 17725 42335
rect 17789 42277 17808 42341
rect 15840 42271 15904 42277
rect 15764 42260 15904 42271
rect 17712 42264 17808 42277
rect 18428 42252 18618 42260
rect 19166 42258 19180 42374
rect 19290 42362 19316 42374
rect 23910 42362 23936 42384
rect 19290 42302 23936 42362
rect 19290 42258 19316 42302
rect 19166 42254 19316 42258
rect 23910 42268 23936 42302
rect 24046 42268 24076 42384
rect 24200 42308 24208 42428
rect 23910 42254 24076 42268
rect 15948 42192 16036 42210
rect 16972 42192 17060 42196
rect 15948 42188 17060 42192
rect 15948 42124 15960 42188
rect 16024 42180 17060 42188
rect 16024 42132 16988 42180
rect 16024 42124 16036 42132
rect 15948 42114 16036 42124
rect 16972 42116 16988 42132
rect 17052 42116 17060 42180
rect 16972 42100 17060 42116
rect 18428 42070 18460 42252
rect 18604 42192 18618 42252
rect 24192 42248 24208 42308
rect 18604 42162 18648 42192
rect 24200 42162 24208 42248
rect 18604 42104 24208 42162
rect 24362 42104 24376 42428
rect 18604 42102 24376 42104
rect 18604 42070 18618 42102
rect 24200 42098 24376 42102
rect 18428 42056 18618 42070
rect 16272 42000 17146 42005
rect 16272 41914 16282 42000
rect 17136 41982 17146 42000
rect 26190 41982 26200 42276
rect 17136 41930 26200 41982
rect 26342 41982 26352 42276
rect 26342 41930 26354 41982
rect 17136 41922 26354 41930
rect 17136 41914 17146 41922
rect 16272 41909 17146 41914
rect 22998 41828 23472 41833
rect 22998 41824 23008 41828
rect 9422 41822 23008 41824
rect 8532 41821 23008 41822
rect 1814 41812 2452 41817
rect 1814 41312 1824 41812
rect 2442 41312 2452 41812
rect 3844 41758 5070 41763
rect 3844 41376 3854 41758
rect 5060 41376 5070 41758
rect 3844 41371 5070 41376
rect 8532 41323 8533 41821
rect 9031 41800 23008 41821
rect 9031 41332 16434 41800
rect 16798 41332 23008 41800
rect 9031 41324 23008 41332
rect 9031 41323 9148 41324
rect 8532 41322 9148 41323
rect 8533 41317 9031 41322
rect 1814 41307 2452 41312
rect 16912 41242 17056 41247
rect 16912 40746 16922 41242
rect 17046 40746 17056 41242
rect 22998 41134 23008 41324
rect 23462 41134 23472 41828
rect 22998 41129 23472 41134
rect 23400 40998 23686 41003
rect 23400 40784 23410 40998
rect 23676 40784 23686 40998
rect 23400 40779 23686 40784
rect 25954 40982 26194 40987
rect 16912 40741 17056 40746
rect 25954 40576 25964 40982
rect 26184 40576 26194 40982
rect 25954 40571 26194 40576
rect 9786 39912 9796 40418
rect 10514 40412 10524 40418
rect 11106 40412 11626 40417
rect 17072 40416 17444 40421
rect 17072 40412 17082 40416
rect 10514 39912 11116 40412
rect 11616 39912 17082 40412
rect 11106 39907 11626 39912
rect 17072 39908 17082 39912
rect 17434 40412 17444 40416
rect 17434 39912 23417 40412
rect 17434 39908 17444 39912
rect 17072 39903 17444 39908
rect 9810 39792 10070 39797
rect 9810 39320 9820 39792
rect 10060 39320 10070 39792
rect 9810 39315 10070 39320
rect 15940 39344 16054 39354
rect 15940 39254 15956 39344
rect 16032 39254 16054 39344
rect 15940 38826 16054 39254
rect 22142 39108 22336 39113
rect 18856 39102 19076 39107
rect 18856 38902 18866 39102
rect 19066 38902 19076 39102
rect 18856 38897 19076 38902
rect 22142 38884 22152 39108
rect 22326 38884 22336 39108
rect 22142 38879 22336 38884
rect 15940 38736 15956 38826
rect 16032 38736 16054 38826
rect 15946 38734 16050 38736
rect 27256 37387 27582 37390
rect 27230 37382 27588 37387
rect 22128 37362 22332 37367
rect 18674 37326 18924 37331
rect 18674 37126 18684 37326
rect 18884 37126 18924 37326
rect 22128 37160 22138 37362
rect 22322 37160 22332 37362
rect 22128 37155 22332 37160
rect 18674 37121 18924 37126
rect 9768 37028 10148 37033
rect 9768 36676 9778 37028
rect 10138 36676 10148 37028
rect 9768 36671 10148 36676
rect 27230 36622 27240 37382
rect 27578 36622 27588 37382
rect 27230 36617 27588 36622
rect 25018 36505 25618 36514
rect 25014 36500 25902 36505
rect 9760 36320 10498 36325
rect 9760 35400 9770 36320
rect 10488 35400 10498 36320
rect 25014 36282 25024 36500
rect 25892 36282 25902 36500
rect 25014 36277 25902 36282
rect 9760 35395 10498 35400
rect 190 34118 200 34990
rect 1668 34898 1678 34990
rect 25018 34898 25618 36277
rect 27256 36125 27582 36617
rect 26520 36120 27608 36125
rect 26520 35632 26530 36120
rect 27598 35632 27608 36120
rect 26520 35627 27608 35632
rect 1668 34298 25636 34898
rect 1668 34118 1678 34298
rect 192 6768 1026 6773
rect 192 6082 202 6768
rect 1016 6082 1026 6768
rect 192 6077 1026 6082
rect 27358 4896 27652 4901
rect 27358 4602 27368 4896
rect 27642 4602 27652 4896
rect 27358 4597 27652 4602
rect 25364 4048 25696 4053
rect 25364 3702 25374 4048
rect 25686 3702 25696 4048
rect 25364 3697 25696 3702
rect 19316 3630 19786 3635
rect 19316 3412 19326 3630
rect 19776 3412 19786 3630
rect 19316 3407 19786 3412
rect 29442 3316 29670 3321
rect 29442 3084 29452 3316
rect 29660 3084 29670 3316
rect 31156 3288 31418 3293
rect 31156 3190 31166 3288
rect 29442 3079 29670 3084
rect 31050 3070 31166 3190
rect 31156 3022 31166 3070
rect 31408 3190 31418 3288
rect 31408 3070 31824 3190
rect 31408 3022 31418 3070
rect 31156 3017 31418 3022
rect 29386 2456 29618 2461
rect 29386 2184 29396 2456
rect 29608 2184 29618 2456
rect 29386 2179 29618 2184
rect 9784 1482 10598 1487
rect 9784 1036 9794 1482
rect 10588 1036 10598 1482
rect 30557 1078 30675 1083
rect 31704 1078 31824 3070
rect 9784 1031 10598 1036
rect 30556 1077 31824 1078
rect 30556 959 30557 1077
rect 30675 959 31824 1077
rect 30556 958 31824 959
rect 30557 953 30675 958
<< via3 >>
rect 13646 44824 14104 44924
rect 16620 44794 16684 44858
rect 14342 44692 14844 44760
rect 796 44518 860 44582
rect 13036 44568 13474 44632
rect 15874 44628 15938 44692
rect 12194 44500 12258 44504
rect 12184 44440 12258 44500
rect 12866 44440 12930 44504
rect 25638 44478 25752 44692
rect 25902 44666 26022 44856
rect 12184 44436 12248 44440
rect 27292 44350 27356 44414
rect 3360 44032 3424 44096
rect 5210 44020 5282 44244
rect 12168 44178 12650 44242
rect 4476 43764 4540 43828
rect 9802 43624 10098 43864
rect 11002 43728 11228 44052
rect 21964 43784 22240 43892
rect 28006 43844 28126 44402
rect 9782 42438 10122 42874
rect 25692 43260 25844 43412
rect 10842 42368 11122 42578
rect 21316 42474 21534 42700
rect 15776 42271 15840 42335
rect 17725 42277 17789 42341
rect 19180 42258 19290 42374
rect 23936 42268 24046 42384
rect 15960 42124 16024 42188
rect 16988 42116 17052 42180
rect 18460 42070 18604 42252
rect 24208 42104 24362 42428
rect 26200 41930 26342 42276
rect 1824 41312 2442 41812
rect 3854 41376 5060 41758
rect 8533 41323 9031 41821
rect 16922 40746 17046 41242
rect 23410 40784 23676 40998
rect 25964 40576 26184 40982
rect 9796 39912 10514 40418
rect 9820 39320 10060 39792
rect 15956 39254 16032 39344
rect 18866 38902 19066 39102
rect 22152 38884 22326 39108
rect 15956 38736 16032 38826
rect 18684 37126 18884 37326
rect 22138 37160 22322 37362
rect 9778 36676 10138 37028
rect 9770 35400 10488 36320
rect 200 34118 1668 34990
rect 202 6082 1016 6768
rect 27368 4602 27642 4896
rect 25374 3702 25686 4048
rect 19326 3412 19776 3630
rect 29452 3084 29660 3316
rect 29396 2184 29608 2456
rect 9794 1036 10588 1482
rect 30557 959 30675 1077
<< metal4 >>
rect 798 44798 858 45152
rect 1534 44798 1594 45152
rect 798 44738 1594 44798
rect 798 44583 858 44738
rect 795 44582 861 44583
rect 795 44518 796 44582
rect 860 44518 861 44582
rect 795 44517 861 44518
rect 200 44094 500 44152
rect 2270 44094 2330 45152
rect 3006 44094 3066 45152
rect 3359 44096 3425 44097
rect 3359 44094 3360 44096
rect 200 44034 3360 44094
rect 200 41824 500 44034
rect 3359 44032 3360 44034
rect 3424 44032 3425 44096
rect 3359 44031 3425 44032
rect 3742 43824 3802 45152
rect 4478 43829 4538 45152
rect 5214 44245 5274 45152
rect 5209 44244 5283 44245
rect 5209 44020 5210 44244
rect 5282 44020 5283 44244
rect 5209 44019 5283 44020
rect 5950 44026 6010 45152
rect 6686 44952 6746 45152
rect 7422 44952 7482 45152
rect 8158 44250 8218 45152
rect 8894 44334 8954 45152
rect 9630 44952 9690 45152
rect 10366 44952 10426 45152
rect 11102 44502 11162 45152
rect 11838 44952 11898 45152
rect 12193 44504 12259 44505
rect 12193 44502 12194 44504
rect 11102 44500 12194 44502
rect 11102 44442 12184 44500
rect 12178 44438 12184 44442
rect 12258 44440 12259 44504
rect 12183 44436 12184 44438
rect 12248 44439 12259 44440
rect 12248 44436 12249 44439
rect 12183 44435 12249 44436
rect 8878 44274 11168 44334
rect 8158 44208 8224 44250
rect 8158 44148 10898 44208
rect 8158 44144 8218 44148
rect 9800 44026 10100 44042
rect 5950 43966 10100 44026
rect 9800 43864 10100 43966
rect 4475 43828 4541 43829
rect 4475 43824 4476 43828
rect 3742 43764 4476 43824
rect 4540 43824 4541 43828
rect 4540 43764 4562 43824
rect 4475 43763 4541 43764
rect 9800 43624 9802 43864
rect 10098 43624 10100 43864
rect 9800 42875 10100 43624
rect 9781 42874 10123 42875
rect 9781 42438 9782 42874
rect 10122 42438 10123 42874
rect 9781 42437 10123 42438
rect 10838 42579 10898 44148
rect 11108 44053 11168 44274
rect 12574 44243 12634 45152
rect 13310 44633 13370 45152
rect 14046 44925 14106 45152
rect 13645 44924 14106 44925
rect 13645 44824 13646 44924
rect 14104 44888 14106 44924
rect 14104 44824 14105 44888
rect 13645 44823 14105 44824
rect 14782 44774 14842 45152
rect 14338 44760 14852 44774
rect 14338 44692 14342 44760
rect 14844 44692 14852 44760
rect 14338 44682 14852 44692
rect 15518 44690 15578 45152
rect 16254 44856 16314 45152
rect 16619 44858 16685 44859
rect 16619 44856 16620 44858
rect 16254 44796 16620 44856
rect 16619 44794 16620 44796
rect 16684 44794 16685 44858
rect 16619 44793 16685 44794
rect 15873 44692 15939 44693
rect 15873 44690 15874 44692
rect 13035 44632 13475 44633
rect 13035 44568 13036 44632
rect 13474 44568 13475 44632
rect 15518 44630 15874 44690
rect 15873 44628 15874 44630
rect 15938 44628 15939 44692
rect 15873 44627 15939 44628
rect 13035 44567 13475 44568
rect 12865 44504 12931 44505
rect 12865 44498 12866 44504
rect 12850 44440 12866 44498
rect 12930 44502 12931 44504
rect 12930 44498 12942 44502
rect 12930 44440 16180 44498
rect 12850 44438 16180 44440
rect 12167 44242 12651 44243
rect 12167 44178 12168 44242
rect 12650 44178 12651 44242
rect 12167 44177 12651 44178
rect 12574 44166 12634 44177
rect 11001 44052 11229 44053
rect 11001 43728 11002 44052
rect 11228 43728 11229 44052
rect 11001 43727 11229 43728
rect 10838 42578 11123 42579
rect 200 41822 8712 41824
rect 200 41821 9032 41822
rect 200 41812 8533 41821
rect 200 41324 1824 41812
rect 200 34991 500 41324
rect 1823 41312 1824 41324
rect 2442 41758 8533 41812
rect 2442 41376 3854 41758
rect 5060 41376 8533 41758
rect 2442 41324 8533 41376
rect 2442 41312 2443 41324
rect 8438 41323 8533 41324
rect 9031 41323 9032 41821
rect 8438 41322 9032 41323
rect 1823 41311 2443 41312
rect 9800 40419 10100 42437
rect 10838 42412 10842 42578
rect 10841 42368 10842 42412
rect 11122 42368 11123 42578
rect 10841 42367 11123 42368
rect 15775 42335 15841 42336
rect 15775 42271 15776 42335
rect 15840 42271 15841 42335
rect 15775 42270 15841 42271
rect 9795 40418 10515 40419
rect 9795 39912 9796 40418
rect 10514 39912 10515 40418
rect 9795 39911 10515 39912
rect 9800 39792 10100 39911
rect 9800 39320 9820 39792
rect 10060 39320 10100 39792
rect 9800 37029 10100 39320
rect 15778 39072 15838 42270
rect 15959 42188 16025 42189
rect 15959 42124 15960 42188
rect 16024 42124 16025 42188
rect 15959 42123 16025 42124
rect 15962 39345 16022 42123
rect 16120 41248 16180 44438
rect 16990 42181 17050 45152
rect 17726 42352 17786 45152
rect 17712 42341 17808 42352
rect 17712 42277 17725 42341
rect 17789 42277 17808 42341
rect 17712 42264 17808 42277
rect 18462 42253 18522 45152
rect 19198 42375 19258 45152
rect 19934 44952 19994 45152
rect 20670 44952 20730 45152
rect 21406 42701 21466 45152
rect 22142 43893 22202 45152
rect 22878 44952 22938 45152
rect 21963 43892 22241 43893
rect 21963 43784 21964 43892
rect 22240 43784 22241 43892
rect 21963 43783 22241 43784
rect 21315 42700 21535 42701
rect 21315 42474 21316 42700
rect 21534 42474 21535 42700
rect 21315 42473 21535 42474
rect 19179 42374 19291 42375
rect 19179 42258 19180 42374
rect 19290 42258 19291 42374
rect 19179 42257 19291 42258
rect 18459 42252 18605 42253
rect 16987 42180 17053 42181
rect 16987 42116 16988 42180
rect 17052 42116 17053 42180
rect 16987 42115 17053 42116
rect 18459 42070 18460 42252
rect 18604 42070 18605 42252
rect 18459 42069 18605 42070
rect 16120 41242 17054 41248
rect 16120 41188 16922 41242
rect 16921 40746 16922 41188
rect 17046 41188 17054 41242
rect 17046 40746 17050 41188
rect 23614 40999 23674 45152
rect 24350 44952 24410 45152
rect 25086 44952 25146 45152
rect 25822 44952 25882 45152
rect 26558 44882 26618 45152
rect 25901 44856 26023 44857
rect 25637 44692 25753 44693
rect 25637 44478 25638 44692
rect 25752 44478 25753 44692
rect 25901 44666 25902 44856
rect 26022 44666 26023 44856
rect 25901 44665 26023 44666
rect 26232 44822 26618 44882
rect 25637 44477 25753 44478
rect 25692 43413 25752 44477
rect 25691 43412 25845 43413
rect 25691 43260 25692 43412
rect 25844 43260 25845 43412
rect 25691 43259 25845 43260
rect 25692 43250 25752 43259
rect 24207 42428 24363 42429
rect 23954 42385 24014 42388
rect 23935 42384 24047 42385
rect 23935 42268 23936 42384
rect 24046 42268 24047 42384
rect 23935 42267 24047 42268
rect 23936 42264 24042 42267
rect 23409 40998 23677 40999
rect 23409 40784 23410 40998
rect 23676 40784 23677 40998
rect 23409 40783 23677 40784
rect 23614 40776 23674 40783
rect 16921 40745 17050 40746
rect 16990 40718 17050 40745
rect 15955 39344 16033 39345
rect 15955 39254 15956 39344
rect 16032 39254 16033 39344
rect 15955 39253 16033 39254
rect 22151 39108 22327 39109
rect 18865 39102 19067 39103
rect 18865 39072 18866 39102
rect 15778 39012 18866 39072
rect 18836 38974 18866 39012
rect 18865 38902 18866 38974
rect 19066 38902 19067 39102
rect 18865 38901 19067 38902
rect 22151 38884 22152 39108
rect 22326 39010 22327 39108
rect 23982 39010 24042 42264
rect 24207 42104 24208 42428
rect 24362 42104 24363 42428
rect 24207 42103 24363 42104
rect 22326 38950 24048 39010
rect 22326 38884 22327 38950
rect 22151 38883 22327 38884
rect 15938 38826 16064 38836
rect 15938 38736 15956 38826
rect 16032 38736 16064 38826
rect 15938 38722 16064 38736
rect 15955 37281 16022 38722
rect 22137 37362 22323 37363
rect 18683 37326 18885 37327
rect 18683 37281 18684 37326
rect 15955 37209 18684 37281
rect 15955 37208 16015 37209
rect 18683 37126 18684 37209
rect 18884 37126 18885 37326
rect 22137 37160 22138 37362
rect 22322 37292 22323 37362
rect 24300 37292 24360 42103
rect 25962 40983 26022 44665
rect 26232 42277 26292 44822
rect 27294 44415 27354 45152
rect 27291 44414 27357 44415
rect 27291 44350 27292 44414
rect 27356 44350 27357 44414
rect 28030 44403 28090 45152
rect 27291 44349 27357 44350
rect 28005 44402 28127 44403
rect 28005 43844 28006 44402
rect 28126 43844 28127 44402
rect 28005 43843 28127 43844
rect 26199 42276 26343 42277
rect 26199 41930 26200 42276
rect 26342 41930 26343 42276
rect 26199 41929 26343 41930
rect 26232 41924 26292 41929
rect 25962 40982 26185 40983
rect 25962 40820 25964 40982
rect 25963 40576 25964 40820
rect 26184 40576 26185 40982
rect 25963 40575 26185 40576
rect 22322 37232 24360 37292
rect 22322 37160 22323 37232
rect 22137 37159 22323 37160
rect 18683 37125 18885 37126
rect 9777 37028 10139 37029
rect 9777 36676 9778 37028
rect 10138 36676 10139 37028
rect 9777 36675 10139 36676
rect 9800 36321 10100 36675
rect 9769 36320 10489 36321
rect 9769 35400 9770 36320
rect 10488 35400 10489 36320
rect 9769 35399 10489 35400
rect 199 34990 1669 34991
rect 199 34118 200 34990
rect 1668 34118 1669 34990
rect 199 34117 1669 34118
rect 200 6769 500 34117
rect 200 6768 1017 6769
rect 200 6082 202 6768
rect 1016 6082 1017 6768
rect 200 6081 1017 6082
rect 200 1000 500 6081
rect 9800 1483 10100 35399
rect 27367 4896 27643 4897
rect 27367 4808 27368 4896
rect 26934 4688 27368 4808
rect 25373 4048 25687 4049
rect 25373 3702 25374 4048
rect 25686 3702 25687 4048
rect 25373 3701 25687 3702
rect 19325 3630 19777 3631
rect 19325 3530 19326 3630
rect 18064 3412 19326 3530
rect 19776 3412 19777 3630
rect 18064 3411 19777 3412
rect 18064 3410 19754 3411
rect 9793 1482 10589 1483
rect 9793 1036 9794 1482
rect 10588 1036 10589 1482
rect 9793 1035 10589 1036
rect 9800 1000 10100 1035
rect 400 0 520 200
rect 4816 0 4936 200
rect 9232 0 9352 200
rect 13648 0 13768 200
rect 18064 0 18184 3410
rect 25452 888 25572 3701
rect 26934 1792 27054 4688
rect 27367 4602 27368 4688
rect 27642 4602 27643 4896
rect 27367 4601 27643 4602
rect 28766 2418 28826 45152
rect 29502 8666 29563 45150
rect 30238 44952 30298 45152
rect 30974 44952 31034 45152
rect 31710 44952 31770 45152
rect 29501 8039 29564 8666
rect 29502 8037 29563 8039
rect 29503 3317 29563 8037
rect 29451 3316 29661 3317
rect 29451 3084 29452 3316
rect 29660 3084 29661 3316
rect 29451 3083 29661 3084
rect 29395 2456 29609 2457
rect 29395 2418 29396 2456
rect 28766 2358 29396 2418
rect 29395 2184 29396 2358
rect 29608 2184 29609 2456
rect 29395 2183 29609 2184
rect 31312 1792 31432 1800
rect 26934 1672 31440 1792
rect 26934 1660 27054 1672
rect 22480 768 25572 888
rect 26896 1077 30676 1078
rect 26896 959 30557 1077
rect 30675 959 30676 1077
rect 26896 958 30676 959
rect 22480 0 22600 768
rect 26896 0 27016 958
rect 31312 0 31432 1672
use cp  cp_0 ~/pll_ssp_submission/Faisal_Tareq_Zayed_AlObaidi/magic
timestamp 1711545388
transform 1 0 24094 0 1 7332
box 3292 -5232 7098 -1340
use Div  Div_0 ~/pll_ssp_submission/Khowla_Alkhulayfi
timestamp 1712557532
transform 1 0 2194 0 -1 42140
box -670 -832 6794 -38
use divi_v1L  divi_v1L_0 ~/pll_ssp_submission/Nawaf/Design_Files/Design_Files/Frequency_Divider
timestamp 1712557532
transform 1 0 980 0 1 40194
box 974 -588 8440 630
use divider  divider_0 ~/pll_ssp_submission/Abdulrahman_Alghamdi/freq_divider
timestamp 1712557532
transform -1 0 23266 0 1 40038
box -200 448 6210 1296
use NFD  NFD_0 ~/pll_ssp_submission/Khalid_Abdulaziz_Mohammed_Al_Zahrani/magic
timestamp 1712557532
transform 0 -1 25184 1 0 36244
box 42 -2334 7908 -1142
use Npfd  Npfd_0 ~/pll_ssp_submission/Baraa_Musa_Abdullah_Al_Harbi/magic
timestamp 1712557532
transform -1 0 23222 0 1 38894
box 1024 -2182 4496 646
use Osc_v3_L  Osc_v3_L_0 ~/pll_ssp_submission/Nawaf/Design_Files/Design_Files/CurrentStarvedOscillator
timestamp 1712227994
transform -1 0 29132 0 1 3170
box 3508 -2212 9578 2934
use pfd_with_buffers  pfd_with_buffers_0 ~/pll_ssp_submission/Abdulrahman_Alghamdi/pfd
timestamp 1712557532
transform -1 0 17586 0 1 43836
box 1572 -1860 6566 514
<< labels >>
flabel metal4 200 1000 500 44152 1 FreeSans 2 0 0 0 VPWR
port 51 nsew power bidirectional
flabel metal4 s 12574 44952 12634 45152 0 FreeSans 480 90 0 0 uo_out[7]
port 50 nsew signal output
flabel metal4 s 13310 44952 13370 45152 0 FreeSans 480 90 0 0 uo_out[6]
port 49 nsew signal output
flabel metal4 s 14046 44952 14106 45152 0 FreeSans 480 90 0 0 uo_out[5]
port 48 nsew signal output
flabel metal4 s 14782 44952 14842 45152 0 FreeSans 480 90 0 0 uo_out[4]
port 47 nsew signal output
flabel metal4 s 15518 44952 15578 45152 0 FreeSans 480 90 0 0 uo_out[3]
port 46 nsew signal output
flabel metal4 s 16254 44952 16314 45152 0 FreeSans 480 90 0 0 uo_out[2]
port 45 nsew signal output
flabel metal4 s 17726 44952 17786 45152 0 FreeSans 480 90 0 0 uo_out[0]
port 43 nsew signal output
flabel metal4 s 6686 44952 6746 45152 0 FreeSans 480 90 0 0 uio_out[7]
port 42 nsew signal output
flabel metal4 s 7422 44952 7482 45152 0 FreeSans 480 90 0 0 uio_out[6]
port 41 nsew signal output
flabel metal4 s 8158 44952 8218 45152 0 FreeSans 480 90 0 0 uio_out[5]
port 40 nsew signal output
flabel metal4 s 8894 44952 8954 45152 0 FreeSans 480 90 0 0 uio_out[4]
port 39 nsew signal output
flabel metal4 s 9630 44952 9690 45152 0 FreeSans 480 90 0 0 uio_out[3]
port 38 nsew signal output
flabel metal4 s 10366 44952 10426 45152 0 FreeSans 480 90 0 0 uio_out[2]
port 37 nsew signal output
flabel metal4 s 11102 44952 11162 45152 0 FreeSans 480 90 0 0 uio_out[1]
port 36 nsew signal output
flabel metal4 s 11838 44952 11898 45152 0 FreeSans 480 90 0 0 uio_out[0]
port 35 nsew signal output
flabel metal4 s 798 44952 858 45152 0 FreeSans 480 90 0 0 uio_oe[7]
port 34 nsew signal output
flabel metal4 s 1534 44952 1594 45152 0 FreeSans 480 90 0 0 uio_oe[6]
port 33 nsew signal output
flabel metal4 s 2270 44952 2330 45152 0 FreeSans 480 90 0 0 uio_oe[5]
port 32 nsew signal output
flabel metal4 s 3006 44952 3066 45152 0 FreeSans 480 90 0 0 uio_oe[4]
port 31 nsew signal output
flabel metal4 s 5214 44952 5274 45152 0 FreeSans 480 90 0 0 uio_oe[1]
port 28 nsew signal output
flabel metal4 s 18462 44952 18522 45152 0 FreeSans 480 90 0 0 uio_in[7]
port 26 nsew signal input
flabel metal4 s 19198 44952 19258 45152 0 FreeSans 480 90 0 0 uio_in[6]
port 25 nsew signal input
flabel metal4 s 19934 44952 19994 45152 0 FreeSans 480 90 0 0 uio_in[5]
port 24 nsew signal input
flabel metal4 s 20670 44952 20730 45152 0 FreeSans 480 90 0 0 uio_in[4]
port 23 nsew signal input
flabel metal4 s 21406 44952 21466 45152 0 FreeSans 480 90 0 0 uio_in[3]
port 22 nsew signal input
flabel metal4 s 22142 44952 22202 45152 0 FreeSans 480 90 0 0 uio_in[2]
port 21 nsew signal input
flabel metal4 s 22878 44952 22938 45152 0 FreeSans 480 90 0 0 uio_in[1]
port 20 nsew signal input
flabel metal4 s 23614 44952 23674 45152 0 FreeSans 480 90 0 0 uio_in[0]
port 19 nsew signal input
flabel metal4 s 24350 44952 24410 45152 0 FreeSans 480 90 0 0 ui_in[7]
port 18 nsew signal input
flabel metal4 s 25086 44952 25146 45152 0 FreeSans 480 90 0 0 ui_in[6]
port 17 nsew signal input
flabel metal4 s 25822 44952 25882 45152 0 FreeSans 480 90 0 0 ui_in[5]
port 16 nsew signal input
flabel metal4 s 26558 44952 26618 45152 0 FreeSans 480 90 0 0 ui_in[4]
port 15 nsew signal input
flabel metal4 s 27294 44952 27354 45152 0 FreeSans 480 90 0 0 ui_in[3]
port 14 nsew signal input
flabel metal4 s 28030 44952 28090 45152 0 FreeSans 480 90 0 0 ui_in[2]
port 13 nsew signal input
flabel metal4 s 28766 44952 28826 45152 0 FreeSans 480 90 0 0 ui_in[1]
port 12 nsew signal input
flabel metal4 s 400 0 520 200 0 FreeSans 960 0 0 0 ua[7]
port 10 nsew signal bidirectional
flabel metal4 s 4816 0 4936 200 0 FreeSans 960 0 0 0 ua[6]
port 9 nsew signal bidirectional
flabel metal4 s 9232 0 9352 200 0 FreeSans 960 0 0 0 ua[5]
port 8 nsew signal bidirectional
flabel metal4 s 13648 0 13768 200 0 FreeSans 960 0 0 0 ua[4]
port 7 nsew signal bidirectional
flabel metal4 s 18064 0 18184 200 0 FreeSans 960 0 0 0 ua[3]
port 6 nsew signal bidirectional
flabel metal4 s 22480 0 22600 200 0 FreeSans 960 0 0 0 ua[2]
port 5 nsew signal bidirectional
flabel metal4 s 26896 0 27016 200 0 FreeSans 960 0 0 0 ua[1]
port 4 nsew signal bidirectional
flabel metal4 s 31312 0 31432 200 0 FreeSans 960 0 0 0 ua[0]
port 3 nsew signal bidirectional
flabel metal4 s 30238 44952 30298 45152 0 FreeSans 480 90 0 0 rst_n
port 2 nsew signal input
flabel metal4 s 31710 44952 31770 45152 0 FreeSans 480 90 0 0 ena
port 1 nsew signal input
flabel metal4 s 30974 44952 31034 45152 0 FreeSans 480 90 0 0 clk
port 0 nsew signal input
flabel metal4 s 16990 44952 17050 45152 0 FreeSans 480 90 0 0 uo_out[1]
port 44 nsew signal output
flabel metal4 s 4478 44952 4538 45152 0 FreeSans 480 90 0 0 uio_oe[2]
port 29 nsew signal output
flabel metal4 s 3742 44952 3802 45152 0 FreeSans 480 90 0 0 uio_oe[3]
port 30 nsew signal output
flabel metal4 s 5950 44952 6010 45152 0 FreeSans 480 90 0 0 uio_oe[0]
port 27 nsew signal output
flabel space 9800 1000 10100 44152 1 FreeSans 2 0 0 0 VGND
port 52 nsew ground bidirectional
flabel metal4 s 29502 44950 29562 45150 0 FreeSans 480 90 0 0 ui_in[0]
port 11 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 32200 45152
<< end >>
