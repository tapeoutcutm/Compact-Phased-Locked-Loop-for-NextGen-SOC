magic
tech sky130A
magscale 1 2
timestamp 1712737205
<< error_p >>
rect -147 681 -89 687
rect -29 681 29 687
rect 89 681 147 687
rect -147 647 -135 681
rect -29 647 -17 681
rect 89 647 101 681
rect -147 641 -89 647
rect -29 641 29 647
rect 89 641 147 647
rect -147 -647 -89 -641
rect -29 -647 29 -641
rect 89 -647 147 -641
rect -147 -681 -135 -647
rect -29 -681 -17 -647
rect 89 -681 101 -647
rect -147 -687 -89 -681
rect -29 -687 29 -681
rect 89 -687 147 -681
<< nwell >>
rect -344 -819 344 819
<< pmos >>
rect -148 -600 -88 600
rect -30 -600 30 600
rect 88 -600 148 600
<< pdiff >>
rect -206 561 -148 600
rect -206 527 -194 561
rect -160 527 -148 561
rect -206 493 -148 527
rect -206 459 -194 493
rect -160 459 -148 493
rect -206 425 -148 459
rect -206 391 -194 425
rect -160 391 -148 425
rect -206 357 -148 391
rect -206 323 -194 357
rect -160 323 -148 357
rect -206 289 -148 323
rect -206 255 -194 289
rect -160 255 -148 289
rect -206 221 -148 255
rect -206 187 -194 221
rect -160 187 -148 221
rect -206 153 -148 187
rect -206 119 -194 153
rect -160 119 -148 153
rect -206 85 -148 119
rect -206 51 -194 85
rect -160 51 -148 85
rect -206 17 -148 51
rect -206 -17 -194 17
rect -160 -17 -148 17
rect -206 -51 -148 -17
rect -206 -85 -194 -51
rect -160 -85 -148 -51
rect -206 -119 -148 -85
rect -206 -153 -194 -119
rect -160 -153 -148 -119
rect -206 -187 -148 -153
rect -206 -221 -194 -187
rect -160 -221 -148 -187
rect -206 -255 -148 -221
rect -206 -289 -194 -255
rect -160 -289 -148 -255
rect -206 -323 -148 -289
rect -206 -357 -194 -323
rect -160 -357 -148 -323
rect -206 -391 -148 -357
rect -206 -425 -194 -391
rect -160 -425 -148 -391
rect -206 -459 -148 -425
rect -206 -493 -194 -459
rect -160 -493 -148 -459
rect -206 -527 -148 -493
rect -206 -561 -194 -527
rect -160 -561 -148 -527
rect -206 -600 -148 -561
rect -88 561 -30 600
rect -88 527 -76 561
rect -42 527 -30 561
rect -88 493 -30 527
rect -88 459 -76 493
rect -42 459 -30 493
rect -88 425 -30 459
rect -88 391 -76 425
rect -42 391 -30 425
rect -88 357 -30 391
rect -88 323 -76 357
rect -42 323 -30 357
rect -88 289 -30 323
rect -88 255 -76 289
rect -42 255 -30 289
rect -88 221 -30 255
rect -88 187 -76 221
rect -42 187 -30 221
rect -88 153 -30 187
rect -88 119 -76 153
rect -42 119 -30 153
rect -88 85 -30 119
rect -88 51 -76 85
rect -42 51 -30 85
rect -88 17 -30 51
rect -88 -17 -76 17
rect -42 -17 -30 17
rect -88 -51 -30 -17
rect -88 -85 -76 -51
rect -42 -85 -30 -51
rect -88 -119 -30 -85
rect -88 -153 -76 -119
rect -42 -153 -30 -119
rect -88 -187 -30 -153
rect -88 -221 -76 -187
rect -42 -221 -30 -187
rect -88 -255 -30 -221
rect -88 -289 -76 -255
rect -42 -289 -30 -255
rect -88 -323 -30 -289
rect -88 -357 -76 -323
rect -42 -357 -30 -323
rect -88 -391 -30 -357
rect -88 -425 -76 -391
rect -42 -425 -30 -391
rect -88 -459 -30 -425
rect -88 -493 -76 -459
rect -42 -493 -30 -459
rect -88 -527 -30 -493
rect -88 -561 -76 -527
rect -42 -561 -30 -527
rect -88 -600 -30 -561
rect 30 561 88 600
rect 30 527 42 561
rect 76 527 88 561
rect 30 493 88 527
rect 30 459 42 493
rect 76 459 88 493
rect 30 425 88 459
rect 30 391 42 425
rect 76 391 88 425
rect 30 357 88 391
rect 30 323 42 357
rect 76 323 88 357
rect 30 289 88 323
rect 30 255 42 289
rect 76 255 88 289
rect 30 221 88 255
rect 30 187 42 221
rect 76 187 88 221
rect 30 153 88 187
rect 30 119 42 153
rect 76 119 88 153
rect 30 85 88 119
rect 30 51 42 85
rect 76 51 88 85
rect 30 17 88 51
rect 30 -17 42 17
rect 76 -17 88 17
rect 30 -51 88 -17
rect 30 -85 42 -51
rect 76 -85 88 -51
rect 30 -119 88 -85
rect 30 -153 42 -119
rect 76 -153 88 -119
rect 30 -187 88 -153
rect 30 -221 42 -187
rect 76 -221 88 -187
rect 30 -255 88 -221
rect 30 -289 42 -255
rect 76 -289 88 -255
rect 30 -323 88 -289
rect 30 -357 42 -323
rect 76 -357 88 -323
rect 30 -391 88 -357
rect 30 -425 42 -391
rect 76 -425 88 -391
rect 30 -459 88 -425
rect 30 -493 42 -459
rect 76 -493 88 -459
rect 30 -527 88 -493
rect 30 -561 42 -527
rect 76 -561 88 -527
rect 30 -600 88 -561
rect 148 561 206 600
rect 148 527 160 561
rect 194 527 206 561
rect 148 493 206 527
rect 148 459 160 493
rect 194 459 206 493
rect 148 425 206 459
rect 148 391 160 425
rect 194 391 206 425
rect 148 357 206 391
rect 148 323 160 357
rect 194 323 206 357
rect 148 289 206 323
rect 148 255 160 289
rect 194 255 206 289
rect 148 221 206 255
rect 148 187 160 221
rect 194 187 206 221
rect 148 153 206 187
rect 148 119 160 153
rect 194 119 206 153
rect 148 85 206 119
rect 148 51 160 85
rect 194 51 206 85
rect 148 17 206 51
rect 148 -17 160 17
rect 194 -17 206 17
rect 148 -51 206 -17
rect 148 -85 160 -51
rect 194 -85 206 -51
rect 148 -119 206 -85
rect 148 -153 160 -119
rect 194 -153 206 -119
rect 148 -187 206 -153
rect 148 -221 160 -187
rect 194 -221 206 -187
rect 148 -255 206 -221
rect 148 -289 160 -255
rect 194 -289 206 -255
rect 148 -323 206 -289
rect 148 -357 160 -323
rect 194 -357 206 -323
rect 148 -391 206 -357
rect 148 -425 160 -391
rect 194 -425 206 -391
rect 148 -459 206 -425
rect 148 -493 160 -459
rect 194 -493 206 -459
rect 148 -527 206 -493
rect 148 -561 160 -527
rect 194 -561 206 -527
rect 148 -600 206 -561
<< pdiffc >>
rect -194 527 -160 561
rect -194 459 -160 493
rect -194 391 -160 425
rect -194 323 -160 357
rect -194 255 -160 289
rect -194 187 -160 221
rect -194 119 -160 153
rect -194 51 -160 85
rect -194 -17 -160 17
rect -194 -85 -160 -51
rect -194 -153 -160 -119
rect -194 -221 -160 -187
rect -194 -289 -160 -255
rect -194 -357 -160 -323
rect -194 -425 -160 -391
rect -194 -493 -160 -459
rect -194 -561 -160 -527
rect -76 527 -42 561
rect -76 459 -42 493
rect -76 391 -42 425
rect -76 323 -42 357
rect -76 255 -42 289
rect -76 187 -42 221
rect -76 119 -42 153
rect -76 51 -42 85
rect -76 -17 -42 17
rect -76 -85 -42 -51
rect -76 -153 -42 -119
rect -76 -221 -42 -187
rect -76 -289 -42 -255
rect -76 -357 -42 -323
rect -76 -425 -42 -391
rect -76 -493 -42 -459
rect -76 -561 -42 -527
rect 42 527 76 561
rect 42 459 76 493
rect 42 391 76 425
rect 42 323 76 357
rect 42 255 76 289
rect 42 187 76 221
rect 42 119 76 153
rect 42 51 76 85
rect 42 -17 76 17
rect 42 -85 76 -51
rect 42 -153 76 -119
rect 42 -221 76 -187
rect 42 -289 76 -255
rect 42 -357 76 -323
rect 42 -425 76 -391
rect 42 -493 76 -459
rect 42 -561 76 -527
rect 160 527 194 561
rect 160 459 194 493
rect 160 391 194 425
rect 160 323 194 357
rect 160 255 194 289
rect 160 187 194 221
rect 160 119 194 153
rect 160 51 194 85
rect 160 -17 194 17
rect 160 -85 194 -51
rect 160 -153 194 -119
rect 160 -221 194 -187
rect 160 -289 194 -255
rect 160 -357 194 -323
rect 160 -425 194 -391
rect 160 -493 194 -459
rect 160 -561 194 -527
<< nsubdiff >>
rect -308 749 -187 783
rect -153 749 -119 783
rect -85 749 -51 783
rect -17 749 17 783
rect 51 749 85 783
rect 119 749 153 783
rect 187 749 308 783
rect -308 663 -274 749
rect 274 663 308 749
rect -308 595 -274 629
rect -308 527 -274 561
rect -308 459 -274 493
rect -308 391 -274 425
rect -308 323 -274 357
rect -308 255 -274 289
rect -308 187 -274 221
rect -308 119 -274 153
rect -308 51 -274 85
rect -308 -17 -274 17
rect -308 -85 -274 -51
rect -308 -153 -274 -119
rect -308 -221 -274 -187
rect -308 -289 -274 -255
rect -308 -357 -274 -323
rect -308 -425 -274 -391
rect -308 -493 -274 -459
rect -308 -561 -274 -527
rect -308 -629 -274 -595
rect 274 595 308 629
rect 274 527 308 561
rect 274 459 308 493
rect 274 391 308 425
rect 274 323 308 357
rect 274 255 308 289
rect 274 187 308 221
rect 274 119 308 153
rect 274 51 308 85
rect 274 -17 308 17
rect 274 -85 308 -51
rect 274 -153 308 -119
rect 274 -221 308 -187
rect 274 -289 308 -255
rect 274 -357 308 -323
rect 274 -425 308 -391
rect 274 -493 308 -459
rect 274 -561 308 -527
rect 274 -629 308 -595
rect -308 -749 -274 -663
rect 274 -749 308 -663
rect -308 -783 -187 -749
rect -153 -783 -119 -749
rect -85 -783 -51 -749
rect -17 -783 17 -749
rect 51 -783 85 -749
rect 119 -783 153 -749
rect 187 -783 308 -749
<< nsubdiffcont >>
rect -187 749 -153 783
rect -119 749 -85 783
rect -51 749 -17 783
rect 17 749 51 783
rect 85 749 119 783
rect 153 749 187 783
rect -308 629 -274 663
rect 274 629 308 663
rect -308 561 -274 595
rect -308 493 -274 527
rect -308 425 -274 459
rect -308 357 -274 391
rect -308 289 -274 323
rect -308 221 -274 255
rect -308 153 -274 187
rect -308 85 -274 119
rect -308 17 -274 51
rect -308 -51 -274 -17
rect -308 -119 -274 -85
rect -308 -187 -274 -153
rect -308 -255 -274 -221
rect -308 -323 -274 -289
rect -308 -391 -274 -357
rect -308 -459 -274 -425
rect -308 -527 -274 -493
rect -308 -595 -274 -561
rect 274 561 308 595
rect 274 493 308 527
rect 274 425 308 459
rect 274 357 308 391
rect 274 289 308 323
rect 274 221 308 255
rect 274 153 308 187
rect 274 85 308 119
rect 274 17 308 51
rect 274 -51 308 -17
rect 274 -119 308 -85
rect 274 -187 308 -153
rect 274 -255 308 -221
rect 274 -323 308 -289
rect 274 -391 308 -357
rect 274 -459 308 -425
rect 274 -527 308 -493
rect 274 -595 308 -561
rect -308 -663 -274 -629
rect 274 -663 308 -629
rect -187 -783 -153 -749
rect -119 -783 -85 -749
rect -51 -783 -17 -749
rect 17 -783 51 -749
rect 85 -783 119 -749
rect 153 -783 187 -749
<< poly >>
rect -151 681 -85 697
rect -151 647 -135 681
rect -101 647 -85 681
rect -151 631 -85 647
rect -33 681 33 697
rect -33 647 -17 681
rect 17 647 33 681
rect -33 631 33 647
rect 85 681 151 697
rect 85 647 101 681
rect 135 647 151 681
rect 85 631 151 647
rect -148 600 -88 631
rect -30 600 30 631
rect 88 600 148 631
rect -148 -631 -88 -600
rect -30 -631 30 -600
rect 88 -631 148 -600
rect -151 -647 -85 -631
rect -151 -681 -135 -647
rect -101 -681 -85 -647
rect -151 -697 -85 -681
rect -33 -647 33 -631
rect -33 -681 -17 -647
rect 17 -681 33 -647
rect -33 -697 33 -681
rect 85 -647 151 -631
rect 85 -681 101 -647
rect 135 -681 151 -647
rect 85 -697 151 -681
<< polycont >>
rect -135 647 -101 681
rect -17 647 17 681
rect 101 647 135 681
rect -135 -681 -101 -647
rect -17 -681 17 -647
rect 101 -681 135 -647
<< locali >>
rect -308 749 -187 783
rect -153 749 -119 783
rect -85 749 -51 783
rect -17 749 17 783
rect 51 749 85 783
rect 119 749 153 783
rect 187 749 308 783
rect -308 663 -274 749
rect -151 647 -135 681
rect -101 647 -85 681
rect -33 647 -17 681
rect 17 647 33 681
rect 85 647 101 681
rect 135 647 151 681
rect 274 663 308 749
rect -308 595 -274 629
rect -308 527 -274 561
rect -308 459 -274 493
rect -308 391 -274 425
rect -308 323 -274 357
rect -308 255 -274 289
rect -308 187 -274 221
rect -308 119 -274 153
rect -308 51 -274 85
rect -308 -17 -274 17
rect -308 -85 -274 -51
rect -308 -153 -274 -119
rect -308 -221 -274 -187
rect -308 -289 -274 -255
rect -308 -357 -274 -323
rect -308 -425 -274 -391
rect -308 -493 -274 -459
rect -308 -561 -274 -527
rect -308 -629 -274 -595
rect -194 561 -160 604
rect -194 493 -160 523
rect -194 425 -160 451
rect -194 357 -160 379
rect -194 289 -160 307
rect -194 221 -160 235
rect -194 153 -160 163
rect -194 85 -160 91
rect -194 17 -160 19
rect -194 -19 -160 -17
rect -194 -91 -160 -85
rect -194 -163 -160 -153
rect -194 -235 -160 -221
rect -194 -307 -160 -289
rect -194 -379 -160 -357
rect -194 -451 -160 -425
rect -194 -523 -160 -493
rect -194 -604 -160 -561
rect -76 561 -42 604
rect -76 493 -42 523
rect -76 425 -42 451
rect -76 357 -42 379
rect -76 289 -42 307
rect -76 221 -42 235
rect -76 153 -42 163
rect -76 85 -42 91
rect -76 17 -42 19
rect -76 -19 -42 -17
rect -76 -91 -42 -85
rect -76 -163 -42 -153
rect -76 -235 -42 -221
rect -76 -307 -42 -289
rect -76 -379 -42 -357
rect -76 -451 -42 -425
rect -76 -523 -42 -493
rect -76 -604 -42 -561
rect 42 561 76 604
rect 42 493 76 523
rect 42 425 76 451
rect 42 357 76 379
rect 42 289 76 307
rect 42 221 76 235
rect 42 153 76 163
rect 42 85 76 91
rect 42 17 76 19
rect 42 -19 76 -17
rect 42 -91 76 -85
rect 42 -163 76 -153
rect 42 -235 76 -221
rect 42 -307 76 -289
rect 42 -379 76 -357
rect 42 -451 76 -425
rect 42 -523 76 -493
rect 42 -604 76 -561
rect 160 561 194 604
rect 160 493 194 523
rect 160 425 194 451
rect 160 357 194 379
rect 160 289 194 307
rect 160 221 194 235
rect 160 153 194 163
rect 160 85 194 91
rect 160 17 194 19
rect 160 -19 194 -17
rect 160 -91 194 -85
rect 160 -163 194 -153
rect 160 -235 194 -221
rect 160 -307 194 -289
rect 160 -379 194 -357
rect 160 -451 194 -425
rect 160 -523 194 -493
rect 160 -604 194 -561
rect 274 595 308 629
rect 274 527 308 561
rect 274 459 308 493
rect 274 391 308 425
rect 274 323 308 357
rect 274 255 308 289
rect 274 187 308 221
rect 274 119 308 153
rect 274 51 308 85
rect 274 -17 308 17
rect 274 -85 308 -51
rect 274 -153 308 -119
rect 274 -221 308 -187
rect 274 -289 308 -255
rect 274 -357 308 -323
rect 274 -425 308 -391
rect 274 -493 308 -459
rect 274 -561 308 -527
rect 274 -629 308 -595
rect -308 -749 -274 -663
rect -151 -681 -135 -647
rect -101 -681 -85 -647
rect -33 -681 -17 -647
rect 17 -681 33 -647
rect 85 -681 101 -647
rect 135 -681 151 -647
rect 274 -749 308 -663
rect -308 -783 -187 -749
rect -153 -783 -119 -749
rect -85 -783 -51 -749
rect -17 -783 17 -749
rect 51 -783 85 -749
rect 119 -783 153 -749
rect 187 -783 308 -749
<< viali >>
rect -135 647 -101 681
rect -17 647 17 681
rect 101 647 135 681
rect -194 527 -160 557
rect -194 523 -160 527
rect -194 459 -160 485
rect -194 451 -160 459
rect -194 391 -160 413
rect -194 379 -160 391
rect -194 323 -160 341
rect -194 307 -160 323
rect -194 255 -160 269
rect -194 235 -160 255
rect -194 187 -160 197
rect -194 163 -160 187
rect -194 119 -160 125
rect -194 91 -160 119
rect -194 51 -160 53
rect -194 19 -160 51
rect -194 -51 -160 -19
rect -194 -53 -160 -51
rect -194 -119 -160 -91
rect -194 -125 -160 -119
rect -194 -187 -160 -163
rect -194 -197 -160 -187
rect -194 -255 -160 -235
rect -194 -269 -160 -255
rect -194 -323 -160 -307
rect -194 -341 -160 -323
rect -194 -391 -160 -379
rect -194 -413 -160 -391
rect -194 -459 -160 -451
rect -194 -485 -160 -459
rect -194 -527 -160 -523
rect -194 -557 -160 -527
rect -76 527 -42 557
rect -76 523 -42 527
rect -76 459 -42 485
rect -76 451 -42 459
rect -76 391 -42 413
rect -76 379 -42 391
rect -76 323 -42 341
rect -76 307 -42 323
rect -76 255 -42 269
rect -76 235 -42 255
rect -76 187 -42 197
rect -76 163 -42 187
rect -76 119 -42 125
rect -76 91 -42 119
rect -76 51 -42 53
rect -76 19 -42 51
rect -76 -51 -42 -19
rect -76 -53 -42 -51
rect -76 -119 -42 -91
rect -76 -125 -42 -119
rect -76 -187 -42 -163
rect -76 -197 -42 -187
rect -76 -255 -42 -235
rect -76 -269 -42 -255
rect -76 -323 -42 -307
rect -76 -341 -42 -323
rect -76 -391 -42 -379
rect -76 -413 -42 -391
rect -76 -459 -42 -451
rect -76 -485 -42 -459
rect -76 -527 -42 -523
rect -76 -557 -42 -527
rect 42 527 76 557
rect 42 523 76 527
rect 42 459 76 485
rect 42 451 76 459
rect 42 391 76 413
rect 42 379 76 391
rect 42 323 76 341
rect 42 307 76 323
rect 42 255 76 269
rect 42 235 76 255
rect 42 187 76 197
rect 42 163 76 187
rect 42 119 76 125
rect 42 91 76 119
rect 42 51 76 53
rect 42 19 76 51
rect 42 -51 76 -19
rect 42 -53 76 -51
rect 42 -119 76 -91
rect 42 -125 76 -119
rect 42 -187 76 -163
rect 42 -197 76 -187
rect 42 -255 76 -235
rect 42 -269 76 -255
rect 42 -323 76 -307
rect 42 -341 76 -323
rect 42 -391 76 -379
rect 42 -413 76 -391
rect 42 -459 76 -451
rect 42 -485 76 -459
rect 42 -527 76 -523
rect 42 -557 76 -527
rect 160 527 194 557
rect 160 523 194 527
rect 160 459 194 485
rect 160 451 194 459
rect 160 391 194 413
rect 160 379 194 391
rect 160 323 194 341
rect 160 307 194 323
rect 160 255 194 269
rect 160 235 194 255
rect 160 187 194 197
rect 160 163 194 187
rect 160 119 194 125
rect 160 91 194 119
rect 160 51 194 53
rect 160 19 194 51
rect 160 -51 194 -19
rect 160 -53 194 -51
rect 160 -119 194 -91
rect 160 -125 194 -119
rect 160 -187 194 -163
rect 160 -197 194 -187
rect 160 -255 194 -235
rect 160 -269 194 -255
rect 160 -323 194 -307
rect 160 -341 194 -323
rect 160 -391 194 -379
rect 160 -413 194 -391
rect 160 -459 194 -451
rect 160 -485 194 -459
rect 160 -527 194 -523
rect 160 -557 194 -527
rect -135 -681 -101 -647
rect -17 -681 17 -647
rect 101 -681 135 -647
<< metal1 >>
rect -147 681 -89 687
rect -147 647 -135 681
rect -101 647 -89 681
rect -147 641 -89 647
rect -29 681 29 687
rect -29 647 -17 681
rect 17 647 29 681
rect -29 641 29 647
rect 89 681 147 687
rect 89 647 101 681
rect 135 647 147 681
rect 89 641 147 647
rect -200 557 -154 600
rect -200 523 -194 557
rect -160 523 -154 557
rect -200 485 -154 523
rect -200 451 -194 485
rect -160 451 -154 485
rect -200 413 -154 451
rect -200 379 -194 413
rect -160 379 -154 413
rect -200 341 -154 379
rect -200 307 -194 341
rect -160 307 -154 341
rect -200 269 -154 307
rect -200 235 -194 269
rect -160 235 -154 269
rect -200 197 -154 235
rect -200 163 -194 197
rect -160 163 -154 197
rect -200 125 -154 163
rect -200 91 -194 125
rect -160 91 -154 125
rect -200 53 -154 91
rect -200 19 -194 53
rect -160 19 -154 53
rect -200 -19 -154 19
rect -200 -53 -194 -19
rect -160 -53 -154 -19
rect -200 -91 -154 -53
rect -200 -125 -194 -91
rect -160 -125 -154 -91
rect -200 -163 -154 -125
rect -200 -197 -194 -163
rect -160 -197 -154 -163
rect -200 -235 -154 -197
rect -200 -269 -194 -235
rect -160 -269 -154 -235
rect -200 -307 -154 -269
rect -200 -341 -194 -307
rect -160 -341 -154 -307
rect -200 -379 -154 -341
rect -200 -413 -194 -379
rect -160 -413 -154 -379
rect -200 -451 -154 -413
rect -200 -485 -194 -451
rect -160 -485 -154 -451
rect -200 -523 -154 -485
rect -200 -557 -194 -523
rect -160 -557 -154 -523
rect -200 -600 -154 -557
rect -82 557 -36 600
rect -82 523 -76 557
rect -42 523 -36 557
rect -82 485 -36 523
rect -82 451 -76 485
rect -42 451 -36 485
rect -82 413 -36 451
rect -82 379 -76 413
rect -42 379 -36 413
rect -82 341 -36 379
rect -82 307 -76 341
rect -42 307 -36 341
rect -82 269 -36 307
rect -82 235 -76 269
rect -42 235 -36 269
rect -82 197 -36 235
rect -82 163 -76 197
rect -42 163 -36 197
rect -82 125 -36 163
rect -82 91 -76 125
rect -42 91 -36 125
rect -82 53 -36 91
rect -82 19 -76 53
rect -42 19 -36 53
rect -82 -19 -36 19
rect -82 -53 -76 -19
rect -42 -53 -36 -19
rect -82 -91 -36 -53
rect -82 -125 -76 -91
rect -42 -125 -36 -91
rect -82 -163 -36 -125
rect -82 -197 -76 -163
rect -42 -197 -36 -163
rect -82 -235 -36 -197
rect -82 -269 -76 -235
rect -42 -269 -36 -235
rect -82 -307 -36 -269
rect -82 -341 -76 -307
rect -42 -341 -36 -307
rect -82 -379 -36 -341
rect -82 -413 -76 -379
rect -42 -413 -36 -379
rect -82 -451 -36 -413
rect -82 -485 -76 -451
rect -42 -485 -36 -451
rect -82 -523 -36 -485
rect -82 -557 -76 -523
rect -42 -557 -36 -523
rect -82 -600 -36 -557
rect 36 557 82 600
rect 36 523 42 557
rect 76 523 82 557
rect 36 485 82 523
rect 36 451 42 485
rect 76 451 82 485
rect 36 413 82 451
rect 36 379 42 413
rect 76 379 82 413
rect 36 341 82 379
rect 36 307 42 341
rect 76 307 82 341
rect 36 269 82 307
rect 36 235 42 269
rect 76 235 82 269
rect 36 197 82 235
rect 36 163 42 197
rect 76 163 82 197
rect 36 125 82 163
rect 36 91 42 125
rect 76 91 82 125
rect 36 53 82 91
rect 36 19 42 53
rect 76 19 82 53
rect 36 -19 82 19
rect 36 -53 42 -19
rect 76 -53 82 -19
rect 36 -91 82 -53
rect 36 -125 42 -91
rect 76 -125 82 -91
rect 36 -163 82 -125
rect 36 -197 42 -163
rect 76 -197 82 -163
rect 36 -235 82 -197
rect 36 -269 42 -235
rect 76 -269 82 -235
rect 36 -307 82 -269
rect 36 -341 42 -307
rect 76 -341 82 -307
rect 36 -379 82 -341
rect 36 -413 42 -379
rect 76 -413 82 -379
rect 36 -451 82 -413
rect 36 -485 42 -451
rect 76 -485 82 -451
rect 36 -523 82 -485
rect 36 -557 42 -523
rect 76 -557 82 -523
rect 36 -600 82 -557
rect 154 557 200 600
rect 154 523 160 557
rect 194 523 200 557
rect 154 485 200 523
rect 154 451 160 485
rect 194 451 200 485
rect 154 413 200 451
rect 154 379 160 413
rect 194 379 200 413
rect 154 341 200 379
rect 154 307 160 341
rect 194 307 200 341
rect 154 269 200 307
rect 154 235 160 269
rect 194 235 200 269
rect 154 197 200 235
rect 154 163 160 197
rect 194 163 200 197
rect 154 125 200 163
rect 154 91 160 125
rect 194 91 200 125
rect 154 53 200 91
rect 154 19 160 53
rect 194 19 200 53
rect 154 -19 200 19
rect 154 -53 160 -19
rect 194 -53 200 -19
rect 154 -91 200 -53
rect 154 -125 160 -91
rect 194 -125 200 -91
rect 154 -163 200 -125
rect 154 -197 160 -163
rect 194 -197 200 -163
rect 154 -235 200 -197
rect 154 -269 160 -235
rect 194 -269 200 -235
rect 154 -307 200 -269
rect 154 -341 160 -307
rect 194 -341 200 -307
rect 154 -379 200 -341
rect 154 -413 160 -379
rect 194 -413 200 -379
rect 154 -451 200 -413
rect 154 -485 160 -451
rect 194 -485 200 -451
rect 154 -523 200 -485
rect 154 -557 160 -523
rect 194 -557 200 -523
rect 154 -600 200 -557
rect -147 -647 -89 -641
rect -147 -681 -135 -647
rect -101 -681 -89 -647
rect -147 -687 -89 -681
rect -29 -647 29 -641
rect -29 -681 -17 -647
rect 17 -681 29 -647
rect -29 -687 29 -681
rect 89 -647 147 -641
rect 89 -681 101 -647
rect 135 -681 147 -647
rect 89 -687 147 -681
<< properties >>
string FIXED_BBOX -291 -766 291 766
<< end >>
