magic
tech sky130A
magscale 1 2
timestamp 1713448658
<< locali >>
rect 10738 29444 11156 29864
<< metal1 >>
rect 8414 44850 8734 44862
rect 8414 44670 8452 44850
rect 8696 44670 8734 44850
rect 9086 44730 9678 44736
rect 9086 44678 9100 44730
rect 9152 44678 9164 44730
rect 9216 44678 9228 44730
rect 9280 44678 9292 44730
rect 9344 44678 9356 44730
rect 9408 44678 9420 44730
rect 9472 44678 9484 44730
rect 9536 44678 9548 44730
rect 9600 44678 9612 44730
rect 9664 44678 9678 44730
rect 9086 44672 9678 44678
rect 8414 44658 8734 44670
rect 1540 44426 1772 44430
rect 1348 44402 1972 44426
rect 1348 44286 1378 44402
rect 1942 44286 1972 44402
rect 1348 44262 1972 44286
rect 1540 42396 1772 44262
rect 8622 44214 8682 44658
rect 9096 44214 9156 44672
rect 27996 44373 28136 44402
rect 10384 44236 12680 44272
rect 10384 44214 12191 44236
rect 10898 44212 12191 44214
rect 12148 44208 12191 44212
rect 12150 44184 12191 44208
rect 12243 44184 12255 44236
rect 12307 44184 12319 44236
rect 12371 44184 12383 44236
rect 12435 44184 12447 44236
rect 12499 44184 12511 44236
rect 12563 44184 12575 44236
rect 12627 44208 12680 44236
rect 12627 44184 12660 44208
rect 12150 44178 12660 44184
rect 6180 43066 6334 43086
rect 6180 42886 6199 43066
rect 6315 42886 6334 43066
rect 6180 42866 6334 42886
rect 8622 42878 8682 44154
rect 9096 43298 9156 44154
rect 9372 43519 9486 43524
rect 9372 43467 9403 43519
rect 9455 43467 9486 43519
rect 9372 43455 9486 43467
rect 9372 43403 9403 43455
rect 9455 43403 9486 43455
rect 9372 43391 9486 43403
rect 9372 43339 9403 43391
rect 9455 43339 9486 43391
rect 9372 43327 9486 43339
rect 8868 43270 9168 43298
rect 8868 43218 8896 43270
rect 8948 43218 8960 43270
rect 9012 43218 9024 43270
rect 9076 43218 9088 43270
rect 9140 43218 9168 43270
rect 8868 43190 9168 43218
rect 9372 43275 9403 43327
rect 9455 43275 9486 43327
rect 9372 43263 9486 43275
rect 9372 43211 9403 43263
rect 9455 43211 9486 43263
rect 9372 43199 9486 43211
rect 9372 43147 9403 43199
rect 9455 43147 9486 43199
rect 9372 43135 9486 43147
rect 9372 43083 9403 43135
rect 9455 43083 9486 43135
rect 9372 43071 9486 43083
rect 9372 43019 9403 43071
rect 9455 43019 9486 43071
rect 9372 43007 9486 43019
rect 9372 42955 9403 43007
rect 9455 42955 9486 43007
rect 9372 42950 9486 42955
rect 8814 42810 9292 42832
rect 8814 42566 8835 42810
rect 9271 42566 9292 42810
rect 8814 42544 9292 42566
rect 1828 41812 2398 42284
rect 1814 41312 1851 41812
rect 2415 41312 2452 41812
rect 4392 41758 4592 41764
rect 3844 41753 5070 41758
rect 3844 41381 3855 41753
rect 5059 41381 5070 41753
rect 3844 41376 5070 41381
rect 4392 40624 4592 41376
rect 9392 41158 9452 42950
rect 6192 41098 9452 41158
rect 6192 40676 6252 41098
rect 10444 40766 10552 44154
rect 10992 44044 11238 44052
rect 10992 43736 11025 44044
rect 11205 43736 11238 44044
rect 15906 43864 22250 43892
rect 15906 43812 21980 43864
rect 22032 43812 22044 43864
rect 22096 43812 22108 43864
rect 22160 43812 22172 43864
rect 22224 43812 22250 43864
rect 27996 43873 28008 44373
rect 28124 43873 28136 44373
rect 27996 43844 28136 43873
rect 15906 43784 22250 43812
rect 10992 43728 11238 43736
rect 15542 43530 15674 43698
rect 15524 43519 15686 43530
rect 15524 42763 15547 43519
rect 15663 42763 15686 43519
rect 25676 43412 25860 43426
rect 25676 43394 26502 43412
rect 25676 43278 25710 43394
rect 25826 43278 26502 43394
rect 25676 43260 26502 43278
rect 25676 43246 25860 43260
rect 15524 42752 15686 42763
rect 10832 42563 11132 42578
rect 10832 42383 10860 42563
rect 11104 42383 11132 42563
rect 10832 42368 11132 42383
rect 8620 40658 10552 40766
rect 1600 40541 1782 40558
rect 1600 39977 1633 40541
rect 1749 40260 1782 40541
rect 11280 40412 11480 42238
rect 15542 41822 15674 42752
rect 21276 42677 21614 42762
rect 21276 42622 21335 42677
rect 15808 42497 21335 42622
rect 21515 42497 21614 42677
rect 15808 42490 21614 42497
rect 21276 42448 21614 42490
rect 22998 41827 23472 41828
rect 15050 41336 15060 41822
rect 15678 41336 15688 41822
rect 16424 41784 16808 41800
rect 16424 41348 16462 41784
rect 16770 41348 16808 41784
rect 15542 41320 15674 41336
rect 16424 41332 16808 41348
rect 1749 40060 2154 40260
rect 1749 39977 1808 40060
rect 1600 39960 1808 39977
rect 1608 39956 1808 39960
rect 11106 39912 11116 40412
rect 11616 39912 11626 40412
rect 4386 39774 10088 39806
rect 4386 39606 9850 39774
rect 9810 39338 9850 39606
rect 10030 39606 10088 39774
rect 16492 39640 16692 41332
rect 16912 41212 17056 41242
rect 16912 40776 16926 41212
rect 17042 40942 17056 41212
rect 22998 41135 23017 41827
rect 23453 41135 23472 41827
rect 25960 41627 26200 41644
rect 25960 41255 25990 41627
rect 26170 41384 26200 41627
rect 26170 41255 26500 41384
rect 25960 41240 26500 41255
rect 25960 41238 26200 41240
rect 22998 41134 23472 41135
rect 17086 40942 17274 40986
rect 17042 40786 17274 40942
rect 23400 40923 23686 40940
rect 17042 40776 17086 40786
rect 16912 40746 17086 40776
rect 16918 40742 17086 40746
rect 23400 40743 23421 40923
rect 23665 40743 23686 40923
rect 23400 40726 23686 40743
rect 17118 40416 17318 40686
rect 17072 40412 17444 40416
rect 17072 39912 17104 40412
rect 17412 39912 17444 40412
rect 17072 39908 17444 39912
rect 10030 39338 10070 39606
rect 16492 39440 21882 39640
rect 9810 39320 10070 39338
rect 18856 39092 19076 39102
rect 18856 38912 18876 39092
rect 19056 38912 19076 39092
rect 18856 38902 19076 38912
rect 22142 39086 22336 39108
rect 22142 38906 22181 39086
rect 22297 38906 22336 39086
rect 22142 38884 22336 38906
rect 27256 38694 27614 38696
rect 27256 37938 27281 38694
rect 27589 37938 27614 38694
rect 27256 37936 27614 37938
rect 25036 37770 25924 37784
rect 25036 37765 26548 37770
rect 25036 37585 25070 37765
rect 25890 37585 26548 37765
rect 28028 37698 28096 43844
rect 26872 37630 28096 37698
rect 28028 37610 28096 37630
rect 25036 37570 26548 37585
rect 25036 37566 25924 37570
rect 22128 37351 22332 37362
rect 18674 37316 18924 37326
rect 18674 37136 18694 37316
rect 18874 37136 18924 37316
rect 22128 37171 22140 37351
rect 22320 37171 22332 37351
rect 22128 37160 22332 37171
rect 18674 37126 18924 37136
rect 9768 37006 10148 37028
rect 9768 36698 9804 37006
rect 10112 36954 10148 37006
rect 10112 36752 19303 36954
rect 10112 36698 10148 36752
rect 9768 36676 10148 36698
rect 9760 36302 10498 36320
rect 9760 35418 9783 36302
rect 10475 36136 10498 36302
rect 10475 36128 26530 36136
rect 10475 36120 27602 36128
rect 10475 36007 27608 36120
rect 10475 35635 26558 36007
rect 27570 35635 27608 36007
rect 10475 35632 27608 35635
rect 10475 35536 26530 35632
rect 10475 35418 10498 35536
rect 9760 35400 10498 35418
rect 28744 35024 28754 35688
rect 28834 35024 28844 35688
rect 28758 33771 28836 35024
rect 29480 35014 29490 35716
rect 29594 35014 29604 35716
rect 8108 30784 8118 31064
rect 9526 31060 9536 31064
rect 15392 31060 15672 31066
rect 9526 30784 15672 31060
rect 9518 30780 15672 30784
rect 192 29784 202 30698
rect 2362 30504 2372 30698
rect 2362 30056 14518 30504
rect 15392 30426 15672 30780
rect 2362 29784 2372 30056
rect 10346 29428 10356 29866
rect 11158 29428 11168 29866
rect 16272 25712 16282 26218
rect 16710 25712 16720 26218
rect 28766 6672 28826 33771
rect 22610 6607 23648 6630
rect 22610 6363 22623 6607
rect 23635 6363 23648 6607
rect 22610 6340 23648 6363
rect 28738 6548 28856 6672
rect 23006 5926 23284 6340
rect 28738 6074 28748 6548
rect 28846 6074 28856 6548
rect 29503 6544 29563 35014
rect 29460 6062 29470 6544
rect 29602 6062 29612 6544
rect 27358 4871 27652 4896
rect 27358 4627 27383 4871
rect 27627 4627 27652 4871
rect 27358 4602 27652 4627
rect 25364 4029 25696 4048
rect 25364 3721 25376 4029
rect 25684 3721 25696 4029
rect 25364 3702 25696 3721
rect 19316 3611 19786 3630
rect 19316 3431 19333 3611
rect 19769 3431 19786 3611
rect 19316 3412 19786 3431
rect 29440 3290 29746 3350
rect 29440 3110 29466 3290
rect 29646 3110 29746 3290
rect 29440 3070 29746 3110
rect 31124 3288 31182 3300
rect 31124 3277 31418 3288
rect 31124 3033 31197 3277
rect 31377 3033 31418 3277
rect 31124 3022 31418 3033
rect 31124 3008 31182 3022
rect 29386 2442 29618 2456
rect 29386 2198 29412 2442
rect 29592 2198 29618 2442
rect 29386 2184 29618 2198
rect 21858 694 22086 1184
rect 21680 668 22192 694
rect 21680 552 21718 668
rect 22154 552 22192 668
rect 21680 526 22192 552
<< via1 >>
rect 8452 44670 8696 44850
rect 9100 44678 9152 44730
rect 9164 44678 9216 44730
rect 9228 44678 9280 44730
rect 9292 44678 9344 44730
rect 9356 44678 9408 44730
rect 9420 44678 9472 44730
rect 9484 44678 9536 44730
rect 9548 44678 9600 44730
rect 9612 44678 9664 44730
rect 1378 44286 1942 44402
rect 12191 44184 12243 44236
rect 12255 44184 12307 44236
rect 12319 44184 12371 44236
rect 12383 44184 12435 44236
rect 12447 44184 12499 44236
rect 12511 44184 12563 44236
rect 12575 44184 12627 44236
rect 6199 42886 6315 43066
rect 9403 43467 9455 43519
rect 9403 43403 9455 43455
rect 9403 43339 9455 43391
rect 8896 43218 8948 43270
rect 8960 43218 9012 43270
rect 9024 43218 9076 43270
rect 9088 43218 9140 43270
rect 9403 43275 9455 43327
rect 9403 43211 9455 43263
rect 9403 43147 9455 43199
rect 9403 43083 9455 43135
rect 9403 43019 9455 43071
rect 9403 42955 9455 43007
rect 8835 42566 9271 42810
rect 1851 41312 2415 41812
rect 3855 41381 5059 41753
rect 11025 43736 11205 44044
rect 21980 43812 22032 43864
rect 22044 43812 22096 43864
rect 22108 43812 22160 43864
rect 22172 43812 22224 43864
rect 28008 43873 28124 44373
rect 15547 42763 15663 43519
rect 25710 43278 25826 43394
rect 10860 42383 11104 42563
rect 1633 39977 1749 40541
rect 21335 42497 21515 42677
rect 15060 41336 15678 41822
rect 16462 41348 16770 41784
rect 11116 39912 11616 40412
rect 9850 39338 10030 39774
rect 16926 40776 17042 41212
rect 23017 41135 23453 41827
rect 25990 41255 26170 41627
rect 23421 40743 23665 40923
rect 17104 39912 17412 40412
rect 18876 38912 19056 39092
rect 22181 38906 22297 39086
rect 27281 37938 27589 38694
rect 25070 37585 25890 37765
rect 18694 37136 18874 37316
rect 22140 37171 22320 37351
rect 9804 36698 10112 37006
rect 9783 35418 10475 36302
rect 26558 35635 27570 36007
rect 28754 35024 28834 35688
rect 29490 35014 29594 35716
rect 8118 30784 9526 31064
rect 202 29784 2362 30698
rect 10356 29428 11158 29866
rect 16282 25712 16710 26218
rect 22623 6363 23635 6607
rect 28748 6074 28846 6548
rect 29470 6062 29602 6544
rect 27383 4627 27627 4871
rect 25376 3721 25684 4029
rect 19333 3431 19769 3611
rect 29466 3110 29646 3290
rect 31197 3033 31377 3277
rect 29412 2198 29592 2442
rect 21718 552 22154 668
<< metal2 >>
rect 8424 44850 8724 44872
rect 8424 44828 8452 44850
rect 8696 44828 8724 44850
rect 8424 44692 8426 44828
rect 8722 44692 8724 44828
rect 8424 44670 8452 44692
rect 8696 44670 8724 44692
rect 8424 44648 8724 44670
rect 9096 44732 9668 44746
rect 9096 44730 9114 44732
rect 9170 44730 9194 44732
rect 9250 44730 9274 44732
rect 9330 44730 9354 44732
rect 9410 44730 9434 44732
rect 9490 44730 9514 44732
rect 9570 44730 9594 44732
rect 9650 44730 9668 44732
rect 9096 44678 9100 44730
rect 9344 44678 9354 44730
rect 9410 44678 9420 44730
rect 9664 44678 9668 44730
rect 9096 44676 9114 44678
rect 9170 44676 9194 44678
rect 9250 44676 9274 44678
rect 9330 44676 9354 44678
rect 9410 44676 9434 44678
rect 9490 44676 9514 44678
rect 9570 44676 9594 44678
rect 9650 44676 9668 44678
rect 9096 44662 9668 44676
rect 9304 44587 10148 44604
rect 9304 44531 9338 44587
rect 9394 44531 9418 44587
rect 9474 44531 9498 44587
rect 9554 44531 9578 44587
rect 9634 44531 9658 44587
rect 9714 44531 9738 44587
rect 9794 44531 9818 44587
rect 9874 44531 9898 44587
rect 9954 44531 9978 44587
rect 10034 44531 10058 44587
rect 10114 44531 10148 44587
rect 9304 44514 10148 44531
rect 1358 44412 1962 44436
rect 1358 44402 1392 44412
rect 1928 44402 1962 44412
rect 1358 44286 1378 44402
rect 1942 44286 1962 44402
rect 1358 44276 1392 44286
rect 1928 44276 1962 44286
rect 1358 44252 1962 44276
rect 9394 44214 9454 44514
rect 28006 44391 28126 44412
rect 28006 44373 28038 44391
rect 28094 44373 28126 44391
rect 12168 44238 12650 44252
rect 12168 44182 12181 44238
rect 12237 44236 12261 44238
rect 12317 44236 12341 44238
rect 12397 44236 12421 44238
rect 12477 44236 12501 44238
rect 12557 44236 12581 44238
rect 12243 44184 12255 44236
rect 12317 44184 12319 44236
rect 12499 44184 12501 44236
rect 12563 44184 12575 44236
rect 12237 44182 12261 44184
rect 12317 44182 12341 44184
rect 12397 44182 12421 44184
rect 12477 44182 12501 44184
rect 12557 44182 12581 44184
rect 12637 44182 12650 44238
rect 12168 44168 12650 44182
rect 9394 43534 9454 44154
rect 11002 44044 11228 44062
rect 11002 44038 11025 44044
rect 11205 44038 11228 44044
rect 11002 43742 11007 44038
rect 11223 43742 11228 44038
rect 21964 43866 22240 43902
rect 21964 43864 21994 43866
rect 22050 43864 22074 43866
rect 22130 43864 22154 43866
rect 22210 43864 22240 43866
rect 21964 43812 21980 43864
rect 22224 43812 22240 43864
rect 28006 43873 28008 44373
rect 28124 43873 28126 44373
rect 28006 43855 28038 43873
rect 28094 43855 28126 43873
rect 28006 43834 28126 43855
rect 21964 43810 21994 43812
rect 22050 43810 22074 43812
rect 22130 43810 22154 43812
rect 22210 43810 22240 43812
rect 21964 43774 22240 43810
rect 11002 43736 11025 43742
rect 11205 43736 11228 43742
rect 11002 43718 11228 43736
rect 9382 43519 9476 43534
rect 9382 43467 9403 43519
rect 9455 43467 9476 43519
rect 9382 43455 9476 43467
rect 9382 43403 9403 43455
rect 9455 43403 9476 43455
rect 9382 43391 9476 43403
rect 9382 43339 9403 43391
rect 9455 43339 9476 43391
rect 9382 43327 9476 43339
rect 8878 43272 9158 43308
rect 8878 43270 8910 43272
rect 8966 43270 8990 43272
rect 9046 43270 9070 43272
rect 9126 43270 9158 43272
rect 8878 43218 8896 43270
rect 9140 43218 9158 43270
rect 8878 43216 8910 43218
rect 8966 43216 8990 43218
rect 9046 43216 9070 43218
rect 9126 43216 9158 43218
rect 8878 43180 9158 43216
rect 9382 43275 9403 43327
rect 9455 43275 9476 43327
rect 9382 43263 9476 43275
rect 9382 43211 9403 43263
rect 9455 43211 9476 43263
rect 9382 43199 9476 43211
rect 9382 43147 9403 43199
rect 9455 43147 9476 43199
rect 9382 43135 9476 43147
rect 6190 43084 6324 43096
rect 6190 43066 6229 43084
rect 6285 43066 6324 43084
rect 6190 42886 6199 43066
rect 6315 42886 6324 43066
rect 9382 43083 9403 43135
rect 9455 43083 9476 43135
rect 9382 43071 9476 43083
rect 9382 43019 9403 43071
rect 9455 43019 9476 43071
rect 9382 43007 9476 43019
rect 9382 42955 9403 43007
rect 9455 42955 9476 43007
rect 9382 42940 9476 42955
rect 15534 43529 15676 43540
rect 6190 42868 6229 42886
rect 6285 42868 6324 42886
rect 6190 42856 6324 42868
rect 9782 42844 10122 42884
rect 8824 42824 9282 42842
rect 9782 42824 9804 42844
rect 8824 42810 9804 42824
rect 8824 42566 8835 42810
rect 9271 42566 9804 42810
rect 8824 42542 9804 42566
rect 8824 42534 9282 42542
rect 9782 42468 9804 42542
rect 10100 42468 10122 42844
rect 15534 42753 15537 43529
rect 15673 42753 15676 43529
rect 25692 43404 25844 43422
rect 25692 43268 25700 43404
rect 25836 43268 25844 43404
rect 25692 43250 25844 43268
rect 15534 42742 15676 42753
rect 21300 42695 21558 42732
rect 9782 42428 10122 42468
rect 10842 42563 11122 42588
rect 10842 42383 10860 42563
rect 11104 42383 11122 42563
rect 21300 42479 21317 42695
rect 21533 42479 21558 42695
rect 21300 42454 21558 42479
rect 10842 42358 11122 42383
rect 16282 41985 17136 42010
rect 16282 41982 16321 41985
rect 1622 41929 16321 41982
rect 16377 41929 16401 41985
rect 16457 41929 16481 41985
rect 16537 41929 16561 41985
rect 16617 41929 16641 41985
rect 16697 41929 16721 41985
rect 16777 41929 16801 41985
rect 16857 41929 16881 41985
rect 16937 41929 16961 41985
rect 17017 41929 17041 41985
rect 17097 41929 17136 41985
rect 1622 41922 17136 41929
rect 1622 40568 1682 41922
rect 16282 41904 17136 41922
rect 15060 41822 15678 41832
rect 1824 41812 2442 41822
rect 1824 41790 1851 41812
rect 2415 41790 2442 41812
rect 1824 41334 1825 41790
rect 2441 41334 2442 41790
rect 3854 41755 5060 41768
rect 3854 41753 3869 41755
rect 5045 41753 5060 41755
rect 3854 41381 3855 41753
rect 5059 41381 5060 41753
rect 3854 41379 3869 41381
rect 5045 41379 5060 41381
rect 3854 41366 5060 41379
rect 1824 41312 1851 41334
rect 2415 41312 2442 41334
rect 23008 41827 23462 41838
rect 15060 41326 15678 41336
rect 16434 41794 16798 41810
rect 16434 41784 16468 41794
rect 16764 41784 16798 41794
rect 16434 41348 16462 41784
rect 16770 41348 16798 41784
rect 16434 41338 16468 41348
rect 16764 41338 16798 41348
rect 16434 41322 16798 41338
rect 1824 41302 2442 41312
rect 16922 41222 17046 41252
rect 16922 41212 16956 41222
rect 17012 41212 17046 41222
rect 16922 40776 16926 41212
rect 17042 40776 17046 41212
rect 23008 41135 23017 41827
rect 23453 41135 23462 41827
rect 25970 41629 26190 41654
rect 25970 41253 25972 41629
rect 26188 41253 26190 41629
rect 25970 41228 26190 41253
rect 23008 41124 23462 41135
rect 16922 40766 16956 40776
rect 17012 40766 17046 40776
rect 16922 40736 17046 40766
rect 23410 40923 23676 40950
rect 23410 40743 23421 40923
rect 23665 40743 23676 40923
rect 23410 40716 23676 40743
rect 1610 40541 1772 40568
rect 1610 39977 1633 40541
rect 1749 39977 1772 40541
rect 1610 39950 1772 39977
rect 11116 40412 11616 40422
rect 11116 39902 11616 39912
rect 17082 40412 17434 40426
rect 17082 39912 17104 40412
rect 17412 39912 17434 40412
rect 17082 39898 17434 39912
rect 9820 39784 10060 39802
rect 9820 39328 9832 39784
rect 10048 39328 10060 39784
rect 9820 39310 10060 39328
rect 18866 39092 19066 39112
rect 18866 38912 18876 39092
rect 19056 38912 19066 39092
rect 18866 38892 19066 38912
rect 22152 39104 22326 39118
rect 22152 38888 22171 39104
rect 22307 38888 22326 39104
rect 22152 38874 22326 38888
rect 27266 38694 27604 38706
rect 27266 37938 27281 38694
rect 27589 37938 27604 38694
rect 27266 37926 27604 37938
rect 25046 37783 25914 37794
rect 25046 37567 25052 37783
rect 25908 37567 25914 37783
rect 25046 37556 25914 37567
rect 22138 37351 22322 37372
rect 18684 37316 18884 37336
rect 18684 37136 18694 37316
rect 18874 37136 18884 37316
rect 22138 37171 22140 37351
rect 22320 37171 22322 37351
rect 22138 37150 22322 37171
rect 18684 37116 18884 37136
rect 9778 37006 10138 37038
rect 9778 36698 9804 37006
rect 10112 36698 10138 37006
rect 9778 36666 10138 36698
rect 9770 36302 10488 36330
rect 9770 36288 9783 36302
rect 10475 36288 10488 36302
rect 9770 35432 9781 36288
rect 10477 35432 10488 36288
rect 26530 36104 27598 36130
rect 26530 35648 26556 36104
rect 27572 35648 27598 36104
rect 29490 35716 29594 35726
rect 26530 35635 26558 35648
rect 27570 35635 27598 35648
rect 26530 35622 27598 35635
rect 28754 35688 28834 35698
rect 9770 35418 9783 35432
rect 10475 35418 10488 35432
rect 9770 35390 10488 35418
rect 28754 35014 28834 35024
rect 29490 35004 29594 35014
rect 8118 31064 9526 31074
rect 8118 30774 9526 30784
rect 202 30698 2362 30708
rect 202 29774 2362 29784
rect 10356 29866 11158 29876
rect 10356 29418 11158 29428
rect 16282 26218 16710 26228
rect 16282 25702 16710 25712
rect 202 6733 1016 6778
rect 202 6117 221 6733
rect 997 6599 1016 6733
rect 22620 6607 23638 6640
rect 22620 6599 22623 6607
rect 997 6363 22623 6599
rect 23635 6599 23638 6607
rect 23635 6596 28415 6599
rect 23635 6363 28426 6596
rect 997 6345 28426 6363
rect 997 6117 1016 6345
rect 22620 6330 23638 6345
rect 202 6072 1016 6117
rect 28036 5612 28426 6345
rect 28748 6548 28846 6558
rect 28748 6064 28846 6074
rect 29470 6544 29602 6554
rect 29470 6052 29602 6062
rect 27368 4871 27642 4906
rect 27368 4627 27383 4871
rect 27627 4627 27642 4871
rect 27368 4592 27642 4627
rect 25374 4029 25686 4058
rect 25374 3721 25376 4029
rect 25684 3721 25686 4029
rect 25374 3692 25686 3721
rect 19326 3629 19776 3640
rect 19326 3611 19363 3629
rect 19739 3611 19776 3629
rect 19326 3431 19333 3611
rect 19769 3431 19776 3611
rect 19326 3413 19363 3431
rect 19739 3413 19776 3431
rect 19326 3402 19776 3413
rect 29452 3308 29660 3326
rect 29452 3290 29488 3308
rect 29624 3290 29660 3308
rect 29452 3110 29466 3290
rect 29646 3110 29660 3290
rect 29452 3092 29488 3110
rect 29624 3092 29660 3110
rect 29452 3074 29660 3092
rect 31166 3277 31408 3298
rect 31166 3263 31197 3277
rect 31377 3263 31408 3277
rect 31166 3047 31179 3263
rect 31395 3047 31408 3263
rect 31166 3033 31197 3047
rect 31377 3033 31408 3047
rect 31166 3012 31408 3033
rect 9794 1447 10588 1492
rect 9794 1071 9803 1447
rect 10579 1071 10588 1447
rect 9794 1026 10588 1071
rect 10332 678 10484 1026
rect 21690 678 22182 704
rect 27588 678 27740 2776
rect 29396 2442 29608 2466
rect 29396 2198 29412 2442
rect 29592 2198 29608 2442
rect 29396 2174 29608 2198
rect 10332 668 27744 678
rect 10332 552 21718 668
rect 22154 552 27744 668
rect 10332 526 27744 552
rect 21690 516 22182 526
<< via2 >>
rect 8426 44692 8452 44828
rect 8452 44692 8696 44828
rect 8696 44692 8722 44828
rect 9114 44730 9170 44732
rect 9194 44730 9250 44732
rect 9274 44730 9330 44732
rect 9354 44730 9410 44732
rect 9434 44730 9490 44732
rect 9514 44730 9570 44732
rect 9594 44730 9650 44732
rect 9114 44678 9152 44730
rect 9152 44678 9164 44730
rect 9164 44678 9170 44730
rect 9194 44678 9216 44730
rect 9216 44678 9228 44730
rect 9228 44678 9250 44730
rect 9274 44678 9280 44730
rect 9280 44678 9292 44730
rect 9292 44678 9330 44730
rect 9354 44678 9356 44730
rect 9356 44678 9408 44730
rect 9408 44678 9410 44730
rect 9434 44678 9472 44730
rect 9472 44678 9484 44730
rect 9484 44678 9490 44730
rect 9514 44678 9536 44730
rect 9536 44678 9548 44730
rect 9548 44678 9570 44730
rect 9594 44678 9600 44730
rect 9600 44678 9612 44730
rect 9612 44678 9650 44730
rect 9114 44676 9170 44678
rect 9194 44676 9250 44678
rect 9274 44676 9330 44678
rect 9354 44676 9410 44678
rect 9434 44676 9490 44678
rect 9514 44676 9570 44678
rect 9594 44676 9650 44678
rect 9338 44531 9394 44587
rect 9418 44531 9474 44587
rect 9498 44531 9554 44587
rect 9578 44531 9634 44587
rect 9658 44531 9714 44587
rect 9738 44531 9794 44587
rect 9818 44531 9874 44587
rect 9898 44531 9954 44587
rect 9978 44531 10034 44587
rect 10058 44531 10114 44587
rect 1392 44402 1928 44412
rect 1392 44286 1928 44402
rect 1392 44276 1928 44286
rect 28038 44373 28094 44391
rect 12181 44236 12237 44238
rect 12261 44236 12317 44238
rect 12341 44236 12397 44238
rect 12421 44236 12477 44238
rect 12501 44236 12557 44238
rect 12581 44236 12637 44238
rect 12181 44184 12191 44236
rect 12191 44184 12237 44236
rect 12261 44184 12307 44236
rect 12307 44184 12317 44236
rect 12341 44184 12371 44236
rect 12371 44184 12383 44236
rect 12383 44184 12397 44236
rect 12421 44184 12435 44236
rect 12435 44184 12447 44236
rect 12447 44184 12477 44236
rect 12501 44184 12511 44236
rect 12511 44184 12557 44236
rect 12581 44184 12627 44236
rect 12627 44184 12637 44236
rect 12181 44182 12237 44184
rect 12261 44182 12317 44184
rect 12341 44182 12397 44184
rect 12421 44182 12477 44184
rect 12501 44182 12557 44184
rect 12581 44182 12637 44184
rect 11007 43742 11025 44038
rect 11025 43742 11205 44038
rect 11205 43742 11223 44038
rect 21994 43864 22050 43866
rect 22074 43864 22130 43866
rect 22154 43864 22210 43866
rect 21994 43812 22032 43864
rect 22032 43812 22044 43864
rect 22044 43812 22050 43864
rect 22074 43812 22096 43864
rect 22096 43812 22108 43864
rect 22108 43812 22130 43864
rect 22154 43812 22160 43864
rect 22160 43812 22172 43864
rect 22172 43812 22210 43864
rect 28038 44335 28094 44373
rect 28038 44255 28094 44311
rect 28038 44175 28094 44231
rect 28038 44095 28094 44151
rect 28038 44015 28094 44071
rect 28038 43935 28094 43991
rect 28038 43873 28094 43911
rect 28038 43855 28094 43873
rect 21994 43810 22050 43812
rect 22074 43810 22130 43812
rect 22154 43810 22210 43812
rect 8910 43270 8966 43272
rect 8990 43270 9046 43272
rect 9070 43270 9126 43272
rect 8910 43218 8948 43270
rect 8948 43218 8960 43270
rect 8960 43218 8966 43270
rect 8990 43218 9012 43270
rect 9012 43218 9024 43270
rect 9024 43218 9046 43270
rect 9070 43218 9076 43270
rect 9076 43218 9088 43270
rect 9088 43218 9126 43270
rect 8910 43216 8966 43218
rect 8990 43216 9046 43218
rect 9070 43216 9126 43218
rect 6229 43066 6285 43084
rect 6229 43028 6285 43066
rect 6229 42948 6285 43004
rect 6229 42886 6285 42924
rect 6229 42868 6285 42886
rect 9804 42468 10100 42844
rect 15537 43519 15673 43529
rect 15537 42763 15547 43519
rect 15547 42763 15663 43519
rect 15663 42763 15673 43519
rect 15537 42753 15673 42763
rect 25700 43394 25836 43404
rect 25700 43278 25710 43394
rect 25710 43278 25826 43394
rect 25826 43278 25836 43394
rect 25700 43268 25836 43278
rect 10874 42405 11090 42541
rect 21317 42677 21533 42695
rect 21317 42497 21335 42677
rect 21335 42497 21515 42677
rect 21515 42497 21533 42677
rect 21317 42479 21533 42497
rect 16321 41929 16377 41985
rect 16401 41929 16457 41985
rect 16481 41929 16537 41985
rect 16561 41929 16617 41985
rect 16641 41929 16697 41985
rect 16721 41929 16777 41985
rect 16801 41929 16857 41985
rect 16881 41929 16937 41985
rect 16961 41929 17017 41985
rect 17041 41929 17097 41985
rect 1825 41334 1851 41790
rect 1851 41334 2415 41790
rect 2415 41334 2441 41790
rect 3869 41753 5045 41755
rect 3869 41381 5045 41753
rect 3869 41379 5045 41381
rect 15060 41336 15678 41822
rect 16468 41784 16764 41794
rect 16468 41348 16764 41784
rect 16468 41338 16764 41348
rect 16956 41212 17012 41222
rect 16956 41166 17012 41212
rect 16956 41086 17012 41142
rect 16956 41006 17012 41062
rect 16956 40926 17012 40982
rect 16956 40846 17012 40902
rect 16956 40776 17012 40822
rect 23047 41173 23423 41789
rect 25972 41627 26188 41629
rect 25972 41255 25990 41627
rect 25990 41255 26170 41627
rect 26170 41255 26188 41627
rect 25972 41253 26188 41255
rect 16956 40766 17012 40776
rect 23435 40765 23651 40901
rect 11138 39934 11594 40390
rect 17110 39934 17406 40390
rect 9832 39774 10048 39784
rect 9832 39338 9850 39774
rect 9850 39338 10030 39774
rect 10030 39338 10048 39774
rect 9832 39328 10048 39338
rect 18898 38934 19034 39070
rect 22171 39086 22307 39104
rect 22171 38906 22181 39086
rect 22181 38906 22297 39086
rect 22297 38906 22307 39086
rect 22171 38888 22307 38906
rect 27287 37968 27583 38664
rect 25052 37765 25908 37783
rect 25052 37585 25070 37765
rect 25070 37585 25890 37765
rect 25890 37585 25908 37765
rect 25052 37567 25908 37585
rect 18716 37158 18852 37294
rect 22162 37193 22298 37329
rect 9810 36704 10106 37000
rect 9781 35432 9783 36288
rect 9783 35432 10475 36288
rect 10475 35432 10477 36288
rect 26556 36007 27572 36104
rect 26556 35648 26558 36007
rect 26558 35648 27570 36007
rect 27570 35648 27572 36007
rect 28754 35024 28834 35688
rect 29490 35014 29594 35716
rect 8118 30784 9526 31064
rect 202 29784 2362 30698
rect 10356 29428 11158 29866
rect 16282 25712 16710 26218
rect 221 6117 997 6733
rect 28748 6074 28846 6548
rect 29470 6062 29602 6544
rect 27397 4641 27613 4857
rect 25382 3727 25678 4023
rect 19363 3611 19739 3629
rect 19363 3431 19739 3611
rect 19363 3413 19739 3431
rect 29488 3290 29624 3308
rect 29488 3110 29624 3290
rect 29488 3092 29624 3110
rect 31179 3047 31197 3263
rect 31197 3047 31377 3263
rect 31377 3047 31395 3263
rect 9803 1071 10579 1447
rect 29434 2212 29570 2428
<< metal3 >>
rect 13636 44906 14114 44924
rect 13636 44874 13683 44906
rect 8412 44842 13683 44874
rect 13747 44842 13763 44906
rect 13827 44842 13843 44906
rect 13907 44842 13923 44906
rect 13987 44842 14003 44906
rect 14067 44842 14114 44906
rect 8412 44828 14114 44842
rect 8412 44814 8426 44828
rect 8414 44692 8426 44814
rect 8722 44824 14114 44828
rect 16620 44858 16684 44864
rect 8722 44814 14110 44824
rect 8722 44692 8734 44814
rect 16684 44833 26032 44856
rect 16684 44796 25930 44833
rect 16620 44788 16684 44794
rect 14322 44758 14858 44784
rect 14322 44752 14361 44758
rect 9076 44732 14361 44752
rect 9076 44692 9114 44732
rect 8414 44653 8734 44692
rect 9086 44676 9114 44692
rect 9170 44676 9194 44732
rect 9250 44676 9274 44732
rect 9330 44676 9354 44732
rect 9410 44676 9434 44732
rect 9490 44676 9514 44732
rect 9570 44676 9594 44732
rect 9650 44694 14361 44732
rect 14425 44694 14441 44758
rect 14505 44694 14521 44758
rect 14585 44694 14601 44758
rect 14665 44694 14681 44758
rect 14745 44694 14761 44758
rect 14825 44694 14858 44758
rect 25892 44769 25930 44796
rect 25994 44769 26032 44833
rect 25892 44753 26032 44769
rect 9650 44692 14858 44694
rect 15874 44692 15938 44698
rect 9650 44676 9678 44692
rect 9086 44667 9678 44676
rect 10148 44612 13063 44632
rect 10092 44599 13063 44612
rect 9294 44587 13063 44599
rect 790 44518 796 44582
rect 860 44518 866 44582
rect 9294 44531 9338 44587
rect 9394 44531 9418 44587
rect 9474 44531 9498 44587
rect 9554 44531 9578 44587
rect 9634 44531 9658 44587
rect 9714 44531 9738 44587
rect 9794 44531 9818 44587
rect 9874 44531 9898 44587
rect 9954 44531 9978 44587
rect 10034 44531 10058 44587
rect 10114 44572 13063 44587
rect 10114 44531 10290 44572
rect 13026 44568 13063 44572
rect 13127 44568 13143 44632
rect 13207 44568 13223 44632
rect 13287 44568 13303 44632
rect 13367 44568 13383 44632
rect 13447 44568 13484 44632
rect 25628 44690 25762 44692
rect 15938 44657 25762 44690
rect 25892 44689 25930 44753
rect 25994 44689 26032 44753
rect 25892 44666 26032 44689
rect 15938 44630 25663 44657
rect 15874 44622 15938 44628
rect 25628 44593 25663 44630
rect 25727 44593 25762 44657
rect 25628 44577 25762 44593
rect 9294 44519 10290 44531
rect 798 43702 858 44518
rect 10092 44512 10290 44519
rect 25628 44513 25663 44577
rect 25727 44513 25762 44577
rect 12140 44442 12150 44506
rect 12400 44502 12410 44506
rect 12834 44502 12844 44506
rect 12400 44442 12844 44502
rect 12834 44438 12844 44442
rect 13140 44438 13150 44506
rect 25628 44478 25762 44513
rect 1348 44412 1972 44431
rect 1332 44352 1392 44412
rect 1348 44276 1392 44352
rect 1928 44370 1972 44412
rect 27222 44414 27378 44426
rect 27222 44370 27292 44414
rect 1928 44350 27292 44370
rect 27356 44350 27378 44414
rect 1928 44310 27378 44350
rect 1928 44276 1972 44310
rect 27222 44306 27378 44310
rect 27996 44395 28136 44407
rect 27996 44331 28034 44395
rect 28098 44331 28136 44395
rect 27996 44315 28136 44331
rect 1348 44257 1972 44276
rect 27996 44251 28034 44315
rect 28098 44251 28136 44315
rect 5200 44180 5214 44244
rect 5278 44180 5292 44244
rect 12158 44242 12660 44247
rect 5200 44164 5292 44180
rect 3360 44096 3424 44102
rect 5200 44100 5214 44164
rect 5278 44100 5292 44164
rect 8104 44142 8114 44214
rect 8480 44154 10898 44214
rect 12158 44178 12177 44242
rect 12241 44178 12257 44242
rect 12321 44178 12337 44242
rect 12401 44178 12417 44242
rect 12481 44178 12497 44242
rect 12561 44178 12577 44242
rect 12641 44178 12660 44242
rect 12158 44173 12660 44178
rect 27996 44235 28136 44251
rect 27996 44171 28034 44235
rect 28098 44171 28136 44235
rect 27996 44155 28136 44171
rect 8480 44142 8490 44154
rect 5200 44094 5292 44100
rect 3424 44084 5292 44094
rect 3424 44034 5214 44084
rect 3360 44026 3424 44032
rect 5200 44020 5214 44034
rect 5278 44020 5292 44084
rect 10822 43976 10832 44154
rect 10898 43976 10908 44154
rect 27996 44091 28034 44155
rect 28098 44091 28136 44155
rect 27996 44075 28136 44091
rect 10992 44042 11238 44057
rect 4470 43764 4476 43828
rect 4540 43826 4546 43828
rect 9790 43826 9800 43872
rect 4540 43766 9800 43826
rect 4540 43764 4546 43766
rect 9790 43702 9800 43766
rect 798 43642 9800 43702
rect 9790 43624 9800 43642
rect 10106 43624 10116 43872
rect 10992 43738 11003 44042
rect 11227 43738 11238 44042
rect 27996 44011 28034 44075
rect 28098 44011 28136 44075
rect 27996 43995 28136 44011
rect 27996 43931 28034 43995
rect 28098 43931 28136 43995
rect 27996 43915 28136 43931
rect 21954 43870 22250 43897
rect 21954 43806 21990 43870
rect 22054 43806 22070 43870
rect 22134 43806 22150 43870
rect 22214 43806 22250 43870
rect 27996 43851 28034 43915
rect 28098 43851 28136 43915
rect 27996 43839 28136 43851
rect 21954 43779 22250 43806
rect 10992 43723 11238 43738
rect 15524 43529 15686 43535
rect 8868 43272 9168 43303
rect 8868 43250 8910 43272
rect 6226 43216 8910 43250
rect 8966 43216 8990 43272
rect 9046 43216 9070 43272
rect 9126 43216 9168 43272
rect 6226 43190 9168 43216
rect 6226 43091 6286 43190
rect 8868 43185 9168 43190
rect 6180 43084 6334 43091
rect 6180 43028 6229 43084
rect 6285 43028 6334 43084
rect 6180 43004 6334 43028
rect 6180 42948 6229 43004
rect 6285 42948 6334 43004
rect 6180 42924 6334 42948
rect 6180 42868 6229 42924
rect 6285 42868 6334 42924
rect 6180 42861 6334 42868
rect 9746 42410 9756 42906
rect 10174 42410 10184 42906
rect 15524 42753 15537 43529
rect 15673 42753 15686 43529
rect 25682 43408 25854 43417
rect 25682 43264 25696 43408
rect 25840 43264 25854 43408
rect 25682 43255 25854 43264
rect 15524 42747 15686 42753
rect 15542 42706 15674 42747
rect 21306 42699 21544 42705
rect 21306 42695 21353 42699
rect 21497 42695 21544 42699
rect 10832 42545 11132 42583
rect 10832 42401 10870 42545
rect 11094 42401 11132 42545
rect 21306 42479 21317 42695
rect 21533 42479 21544 42695
rect 21306 42475 21353 42479
rect 21497 42475 21544 42479
rect 21306 42469 21544 42475
rect 10832 42363 11132 42401
rect 19166 42362 19316 42384
rect 23910 42362 24076 42398
rect 19166 42358 24076 42362
rect 15764 42337 15904 42352
rect 17712 42341 17808 42352
rect 17712 42337 17725 42341
rect 15764 42335 17725 42337
rect 15764 42271 15776 42335
rect 15840 42277 17725 42335
rect 17789 42277 17808 42341
rect 15840 42271 15904 42277
rect 15764 42260 15904 42271
rect 17712 42264 17808 42277
rect 19166 42348 23959 42358
rect 19166 42284 19203 42348
rect 19267 42302 23959 42348
rect 19267 42284 19316 42302
rect 18428 42233 18618 42260
rect 19166 42254 19316 42284
rect 23910 42294 23959 42302
rect 24023 42294 24076 42358
rect 23910 42254 24076 42294
rect 26190 42255 26352 42276
rect 15948 42192 16036 42210
rect 16972 42192 17060 42196
rect 15948 42188 17060 42192
rect 15948 42124 15960 42188
rect 16024 42180 17060 42188
rect 16024 42132 16988 42180
rect 16024 42124 16036 42132
rect 15948 42114 16036 42124
rect 16972 42116 16988 42132
rect 17052 42116 17060 42180
rect 16972 42100 17060 42116
rect 18428 42089 18460 42233
rect 18604 42192 18618 42233
rect 18604 42162 18648 42192
rect 26190 42191 26239 42255
rect 26303 42191 26352 42255
rect 26190 42175 26352 42191
rect 24178 42162 24410 42166
rect 18604 42146 24410 42162
rect 18604 42102 24222 42146
rect 18604 42089 18618 42102
rect 18428 42056 18618 42089
rect 24178 42082 24222 42102
rect 24286 42082 24302 42146
rect 24366 42082 24410 42146
rect 24178 42062 24410 42082
rect 26190 42111 26239 42175
rect 26303 42111 26352 42175
rect 26190 42095 26352 42111
rect 26190 42031 26239 42095
rect 26303 42031 26352 42095
rect 26190 42015 26352 42031
rect 16272 41985 17146 42005
rect 16272 41929 16321 41985
rect 16377 41929 16401 41985
rect 16457 41929 16481 41985
rect 16537 41929 16561 41985
rect 16617 41929 16641 41985
rect 16697 41929 16721 41985
rect 16777 41929 16801 41985
rect 16857 41929 16881 41985
rect 16937 41929 16961 41985
rect 17017 41929 17041 41985
rect 17097 41982 17146 41985
rect 26190 41982 26239 42015
rect 17097 41951 26239 41982
rect 26303 41982 26352 42015
rect 26303 41951 26354 41982
rect 17097 41929 26354 41951
rect 16272 41922 26354 41929
rect 16272 41909 17146 41922
rect 1798 41288 1808 41838
rect 2480 41288 2490 41838
rect 8533 41824 9031 41827
rect 9798 41824 10102 41832
rect 15050 41824 15688 41827
rect 22998 41824 23472 41833
rect 3844 41755 5070 41763
rect 3844 41719 3869 41755
rect 5045 41719 5070 41755
rect 3844 41415 3865 41719
rect 5049 41415 5070 41719
rect 3844 41379 3869 41415
rect 5045 41379 5070 41415
rect 3844 41371 5070 41379
rect 8524 41324 8530 41824
rect 9030 41822 23472 41824
rect 9030 41336 15060 41822
rect 15678 41794 23472 41822
rect 15678 41338 16468 41794
rect 16764 41789 23472 41794
rect 16764 41338 23047 41789
rect 15678 41336 23047 41338
rect 9030 41324 23047 41336
rect 8532 41322 9148 41324
rect 8533 41317 9031 41322
rect 9798 41314 10102 41324
rect 16912 41226 17056 41247
rect 16912 41162 16952 41226
rect 17016 41162 17056 41226
rect 16912 41146 17056 41162
rect 16912 41082 16952 41146
rect 17016 41082 17056 41146
rect 22998 41173 23047 41324
rect 23423 41173 23472 41789
rect 25960 41633 26200 41649
rect 25960 41629 26008 41633
rect 26152 41629 26200 41633
rect 25960 41253 25972 41629
rect 26188 41253 26200 41629
rect 25960 41249 26008 41253
rect 26152 41249 26200 41253
rect 25960 41233 26200 41249
rect 22998 41129 23472 41173
rect 16912 41066 17056 41082
rect 16912 41002 16952 41066
rect 17016 41002 17056 41066
rect 16912 40986 17056 41002
rect 16912 40922 16952 40986
rect 17016 40922 17056 40986
rect 16912 40906 17056 40922
rect 16912 40842 16952 40906
rect 17016 40842 17056 40906
rect 16912 40826 17056 40842
rect 16912 40762 16952 40826
rect 17016 40762 17056 40826
rect 16912 40741 17056 40762
rect 23400 40905 23686 40945
rect 23400 40761 23431 40905
rect 23655 40761 23686 40905
rect 23400 40721 23686 40761
rect 9786 40412 10524 40418
rect 11106 40412 11626 40417
rect 17072 40412 17444 40421
rect 9786 40397 17472 40412
rect 9786 39933 10100 40397
rect 10507 40390 17472 40397
rect 10507 39934 11138 40390
rect 11594 39934 17110 40390
rect 17406 39934 17472 40390
rect 10507 39933 17472 39934
rect 9786 39912 17472 39933
rect 11106 39907 11626 39912
rect 17072 39903 17444 39912
rect 9810 39784 10070 39797
rect 9810 39328 9832 39784
rect 10048 39328 10070 39784
rect 9810 39315 10070 39328
rect 15940 39331 16054 39354
rect 15940 39267 15962 39331
rect 16026 39267 16054 39331
rect 15940 38813 16054 39267
rect 22142 39108 22336 39113
rect 18856 39074 19076 39107
rect 18856 38930 18894 39074
rect 19038 38930 19076 39074
rect 18856 38897 19076 38930
rect 22142 38884 22167 39108
rect 22311 38884 22336 39108
rect 22142 38879 22336 38884
rect 15940 38749 15962 38813
rect 16026 38749 16054 38813
rect 15940 38736 16054 38749
rect 15946 38734 16050 38736
rect 27282 38701 27608 38704
rect 27256 38664 27614 38701
rect 27256 37968 27287 38664
rect 27583 37968 27614 38664
rect 27256 37931 27614 37968
rect 27256 37896 27608 37931
rect 25018 37798 25618 37834
rect 25018 37789 25640 37798
rect 25018 37783 25924 37789
rect 25018 37567 25052 37783
rect 25908 37567 25924 37783
rect 25018 37561 25924 37567
rect 25018 37522 25640 37561
rect 22128 37333 22332 37367
rect 18674 37298 18924 37331
rect 18674 37154 18712 37298
rect 18856 37154 18924 37298
rect 22128 37189 22158 37333
rect 22302 37189 22332 37333
rect 22128 37155 22332 37189
rect 18674 37121 18924 37154
rect 9744 36664 9754 37054
rect 10188 36664 10198 37054
rect 9760 36292 10498 36325
rect 9760 36288 10100 36292
rect 9760 35432 9781 36288
rect 9760 35428 10100 35432
rect 10481 35428 10498 36292
rect 9760 35395 10498 35428
rect 190 34986 1678 34990
rect 190 34122 222 34986
rect 1646 34898 1678 34986
rect 25018 34898 25618 37522
rect 27256 36125 27582 37896
rect 26520 36104 27608 36125
rect 26520 35648 26556 36104
rect 27572 35648 27608 36104
rect 29480 35716 29604 35721
rect 26520 35627 27608 35648
rect 28744 35688 28844 35693
rect 28744 35024 28754 35688
rect 28834 35024 28844 35688
rect 28744 35019 28844 35024
rect 29480 35014 29490 35716
rect 29594 35014 29604 35716
rect 29480 35009 29604 35014
rect 1646 34298 25636 34898
rect 1646 34122 1678 34298
rect 190 34118 1678 34122
rect 7309 31767 16772 32089
rect 192 30698 2372 30703
rect 192 29784 202 30698
rect 2362 29784 2372 30698
rect 192 29779 2372 29784
rect 192 6737 1026 6773
rect 192 6113 217 6737
rect 1001 6113 1026 6737
rect 192 6077 1026 6113
rect 7309 1881 7631 31767
rect 8148 31069 8428 31070
rect 8108 31064 9536 31069
rect 8108 30784 8118 31064
rect 9526 30784 9536 31064
rect 8108 30779 9536 30784
rect 8148 5766 8428 30779
rect 16450 30717 16772 31767
rect 10346 29866 11168 29871
rect 10346 29428 10356 29866
rect 11158 29428 11168 29866
rect 10346 29423 11168 29428
rect 16272 26218 16720 26223
rect 16272 25712 16282 26218
rect 16710 25712 16720 26218
rect 16272 25707 16720 25712
rect 28738 6548 28856 6553
rect 28738 6074 28748 6548
rect 28846 6074 28856 6548
rect 28738 6069 28856 6074
rect 29460 6544 29612 6549
rect 29460 6062 29470 6544
rect 29602 6062 29612 6544
rect 29460 6057 29612 6062
rect 8148 5444 13851 5766
rect 8148 5406 8428 5444
rect 13529 2792 13851 5444
rect 27358 4861 27652 4901
rect 27358 4637 27393 4861
rect 27617 4637 27652 4861
rect 27358 4597 27652 4637
rect 25364 4027 25696 4053
rect 25364 3723 25378 4027
rect 25682 3723 25696 4027
rect 25364 3697 25696 3723
rect 19316 3629 19786 3635
rect 19316 3593 19363 3629
rect 19739 3593 19786 3629
rect 19316 3449 19359 3593
rect 19743 3449 19786 3593
rect 19316 3413 19363 3449
rect 19739 3413 19786 3449
rect 19316 3407 19786 3413
rect 29442 3312 29670 3321
rect 29442 3088 29484 3312
rect 29628 3088 29670 3312
rect 31156 3263 31418 3293
rect 31156 3190 31179 3263
rect 29442 3079 29670 3088
rect 31050 3070 31179 3190
rect 31156 3047 31179 3070
rect 31395 3190 31418 3263
rect 31395 3070 31824 3190
rect 31395 3047 31418 3070
rect 31156 3017 31418 3047
rect 8156 1881 8166 1900
rect 7309 1559 8166 1881
rect 8156 1554 8166 1559
rect 9398 1554 9408 1900
rect 9784 1451 10598 1487
rect 9784 1447 10100 1451
rect 9784 1071 9803 1447
rect 9784 1067 10100 1071
rect 10583 1067 10598 1451
rect 9784 1031 10598 1067
rect 13514 1062 13524 2792
rect 13892 1062 13902 2792
rect 29386 2432 29618 2461
rect 29386 2208 29430 2432
rect 29574 2208 29618 2432
rect 29386 2179 29618 2208
rect 30557 1078 30675 1083
rect 31704 1078 31824 3070
rect 13529 1049 13851 1062
rect 30556 1050 31824 1078
rect 30556 986 30584 1050
rect 30648 986 31824 1050
rect 30556 958 31824 986
rect 30557 953 30675 958
<< via3 >>
rect 13683 44842 13747 44906
rect 13763 44842 13827 44906
rect 13843 44842 13907 44906
rect 13923 44842 13987 44906
rect 14003 44842 14067 44906
rect 16620 44794 16684 44858
rect 14361 44694 14425 44758
rect 14441 44694 14505 44758
rect 14521 44694 14585 44758
rect 14601 44694 14665 44758
rect 14681 44694 14745 44758
rect 14761 44694 14825 44758
rect 25930 44769 25994 44833
rect 796 44518 860 44582
rect 13063 44568 13127 44632
rect 13143 44568 13207 44632
rect 13223 44568 13287 44632
rect 13303 44568 13367 44632
rect 13383 44568 13447 44632
rect 15874 44628 15938 44692
rect 25930 44689 25994 44753
rect 25663 44593 25727 44657
rect 25663 44513 25727 44577
rect 12150 44442 12400 44506
rect 12844 44438 13140 44506
rect 27292 44350 27356 44414
rect 28034 44391 28098 44395
rect 28034 44335 28038 44391
rect 28038 44335 28094 44391
rect 28094 44335 28098 44391
rect 28034 44331 28098 44335
rect 28034 44311 28098 44315
rect 28034 44255 28038 44311
rect 28038 44255 28094 44311
rect 28094 44255 28098 44311
rect 28034 44251 28098 44255
rect 5214 44180 5278 44244
rect 3360 44032 3424 44096
rect 5214 44100 5278 44164
rect 8114 44142 8480 44214
rect 12177 44238 12241 44242
rect 12177 44182 12181 44238
rect 12181 44182 12237 44238
rect 12237 44182 12241 44238
rect 12177 44178 12241 44182
rect 12257 44238 12321 44242
rect 12257 44182 12261 44238
rect 12261 44182 12317 44238
rect 12317 44182 12321 44238
rect 12257 44178 12321 44182
rect 12337 44238 12401 44242
rect 12337 44182 12341 44238
rect 12341 44182 12397 44238
rect 12397 44182 12401 44238
rect 12337 44178 12401 44182
rect 12417 44238 12481 44242
rect 12417 44182 12421 44238
rect 12421 44182 12477 44238
rect 12477 44182 12481 44238
rect 12417 44178 12481 44182
rect 12497 44238 12561 44242
rect 12497 44182 12501 44238
rect 12501 44182 12557 44238
rect 12557 44182 12561 44238
rect 12497 44178 12561 44182
rect 12577 44238 12641 44242
rect 12577 44182 12581 44238
rect 12581 44182 12637 44238
rect 12637 44182 12641 44238
rect 12577 44178 12641 44182
rect 28034 44231 28098 44235
rect 28034 44175 28038 44231
rect 28038 44175 28094 44231
rect 28094 44175 28098 44231
rect 28034 44171 28098 44175
rect 5214 44020 5278 44084
rect 10832 43976 10898 44154
rect 28034 44151 28098 44155
rect 28034 44095 28038 44151
rect 28038 44095 28094 44151
rect 28094 44095 28098 44151
rect 28034 44091 28098 44095
rect 4476 43764 4540 43828
rect 9800 43624 10106 43872
rect 11003 44038 11227 44042
rect 11003 43742 11007 44038
rect 11007 43742 11223 44038
rect 11223 43742 11227 44038
rect 11003 43738 11227 43742
rect 28034 44071 28098 44075
rect 28034 44015 28038 44071
rect 28038 44015 28094 44071
rect 28094 44015 28098 44071
rect 28034 44011 28098 44015
rect 28034 43991 28098 43995
rect 28034 43935 28038 43991
rect 28038 43935 28094 43991
rect 28094 43935 28098 43991
rect 28034 43931 28098 43935
rect 21990 43866 22054 43870
rect 21990 43810 21994 43866
rect 21994 43810 22050 43866
rect 22050 43810 22054 43866
rect 21990 43806 22054 43810
rect 22070 43866 22134 43870
rect 22070 43810 22074 43866
rect 22074 43810 22130 43866
rect 22130 43810 22134 43866
rect 22070 43806 22134 43810
rect 22150 43866 22214 43870
rect 22150 43810 22154 43866
rect 22154 43810 22210 43866
rect 22210 43810 22214 43866
rect 22150 43806 22214 43810
rect 28034 43911 28098 43915
rect 28034 43855 28038 43911
rect 28038 43855 28094 43911
rect 28094 43855 28098 43911
rect 28034 43851 28098 43855
rect 9756 42844 10174 42906
rect 9756 42468 9804 42844
rect 9804 42468 10100 42844
rect 10100 42468 10174 42844
rect 9756 42410 10174 42468
rect 25696 43404 25840 43408
rect 25696 43268 25700 43404
rect 25700 43268 25836 43404
rect 25836 43268 25840 43404
rect 25696 43264 25840 43268
rect 21353 42695 21497 42699
rect 10870 42541 11094 42545
rect 10870 42405 10874 42541
rect 10874 42405 11090 42541
rect 11090 42405 11094 42541
rect 10870 42401 11094 42405
rect 21353 42479 21497 42695
rect 21353 42475 21497 42479
rect 15776 42271 15840 42335
rect 17725 42277 17789 42341
rect 19203 42284 19267 42348
rect 23959 42294 24023 42358
rect 15960 42124 16024 42188
rect 16988 42116 17052 42180
rect 18460 42089 18604 42233
rect 26239 42191 26303 42255
rect 24222 42082 24286 42146
rect 24302 42082 24366 42146
rect 26239 42111 26303 42175
rect 26239 42031 26303 42095
rect 26239 41951 26303 42015
rect 1808 41790 2480 41838
rect 1808 41334 1825 41790
rect 1825 41334 2441 41790
rect 2441 41334 2480 41790
rect 1808 41288 2480 41334
rect 3865 41415 3869 41719
rect 3869 41415 5045 41719
rect 5045 41415 5049 41719
rect 8530 41324 9030 41824
rect 15060 41336 15678 41822
rect 16952 41222 17016 41226
rect 16952 41166 16956 41222
rect 16956 41166 17012 41222
rect 17012 41166 17016 41222
rect 16952 41162 17016 41166
rect 16952 41142 17016 41146
rect 16952 41086 16956 41142
rect 16956 41086 17012 41142
rect 17012 41086 17016 41142
rect 16952 41082 17016 41086
rect 26008 41629 26152 41633
rect 26008 41253 26152 41629
rect 26008 41249 26152 41253
rect 16952 41062 17016 41066
rect 16952 41006 16956 41062
rect 16956 41006 17012 41062
rect 17012 41006 17016 41062
rect 16952 41002 17016 41006
rect 16952 40982 17016 40986
rect 16952 40926 16956 40982
rect 16956 40926 17012 40982
rect 17012 40926 17016 40982
rect 16952 40922 17016 40926
rect 16952 40902 17016 40906
rect 16952 40846 16956 40902
rect 16956 40846 17012 40902
rect 17012 40846 17016 40902
rect 16952 40842 17016 40846
rect 16952 40822 17016 40826
rect 16952 40766 16956 40822
rect 16956 40766 17012 40822
rect 17012 40766 17016 40822
rect 16952 40762 17016 40766
rect 23431 40901 23655 40905
rect 23431 40765 23435 40901
rect 23435 40765 23651 40901
rect 23651 40765 23655 40901
rect 23431 40761 23655 40765
rect 10100 39933 10507 40397
rect 15962 39267 16026 39331
rect 18894 39070 19038 39074
rect 18894 38934 18898 39070
rect 18898 38934 19034 39070
rect 19034 38934 19038 39070
rect 18894 38930 19038 38934
rect 22167 39104 22311 39108
rect 22167 38888 22171 39104
rect 22171 38888 22307 39104
rect 22307 38888 22311 39104
rect 22167 38884 22311 38888
rect 15962 38749 16026 38813
rect 18712 37294 18856 37298
rect 18712 37158 18716 37294
rect 18716 37158 18852 37294
rect 18852 37158 18856 37294
rect 18712 37154 18856 37158
rect 22158 37329 22302 37333
rect 22158 37193 22162 37329
rect 22162 37193 22298 37329
rect 22298 37193 22302 37329
rect 22158 37189 22302 37193
rect 9754 37000 10188 37054
rect 9754 36704 9810 37000
rect 9810 36704 10106 37000
rect 10106 36704 10188 37000
rect 9754 36664 10188 36704
rect 10100 36288 10481 36292
rect 10100 35432 10477 36288
rect 10477 35432 10481 36288
rect 10100 35428 10481 35432
rect 222 34122 1646 34986
rect 28754 35024 28834 35688
rect 29490 35014 29594 35716
rect 202 29784 2362 30698
rect 217 6733 1001 6737
rect 217 6117 221 6733
rect 221 6117 997 6733
rect 997 6117 1001 6733
rect 217 6113 1001 6117
rect 10356 29428 11158 29866
rect 16282 25712 16710 26218
rect 28748 6074 28846 6548
rect 29470 6062 29602 6544
rect 27393 4857 27617 4861
rect 27393 4641 27397 4857
rect 27397 4641 27613 4857
rect 27613 4641 27617 4857
rect 27393 4637 27617 4641
rect 25378 4023 25682 4027
rect 25378 3727 25382 4023
rect 25382 3727 25678 4023
rect 25678 3727 25682 4023
rect 25378 3723 25682 3727
rect 19359 3449 19363 3593
rect 19363 3449 19739 3593
rect 19739 3449 19743 3593
rect 29484 3308 29628 3312
rect 29484 3092 29488 3308
rect 29488 3092 29624 3308
rect 29624 3092 29628 3308
rect 29484 3088 29628 3092
rect 8166 1554 9398 1900
rect 10100 1447 10583 1451
rect 10100 1071 10579 1447
rect 10579 1071 10583 1447
rect 10100 1067 10583 1071
rect 13524 1062 13892 2792
rect 29430 2428 29574 2432
rect 29430 2212 29434 2428
rect 29434 2212 29570 2428
rect 29570 2212 29574 2428
rect 29430 2208 29574 2212
rect 30584 986 30648 1050
<< metal4 >>
rect 798 44798 858 45152
rect 1534 44798 1594 45152
rect 798 44738 1594 44798
rect 798 44583 858 44738
rect 795 44582 861 44583
rect 795 44518 796 44582
rect 860 44518 861 44582
rect 795 44517 861 44518
rect 200 44094 500 44152
rect 2270 44094 2330 45152
rect 3006 44094 3066 45152
rect 3359 44096 3425 44097
rect 3359 44094 3360 44096
rect 200 44034 3360 44094
rect 200 41824 500 44034
rect 3359 44032 3360 44034
rect 3424 44032 3425 44096
rect 3359 44031 3425 44032
rect 3742 43824 3802 45152
rect 4478 43829 4538 45152
rect 5214 44245 5274 45152
rect 5209 44244 5283 44245
rect 5209 44180 5214 44244
rect 5278 44180 5283 44244
rect 5209 44164 5283 44180
rect 5209 44100 5214 44164
rect 5278 44100 5283 44164
rect 5209 44084 5283 44100
rect 5209 44020 5214 44084
rect 5278 44020 5283 44084
rect 5209 44019 5283 44020
rect 5950 44026 6010 45152
rect 6686 44952 6746 45152
rect 7422 44952 7482 45152
rect 8158 44250 8218 45152
rect 8894 44334 8954 45152
rect 9630 44952 9690 45152
rect 10366 44952 10426 45152
rect 11102 44502 11162 45152
rect 11838 44952 11898 45152
rect 12149 44506 12401 44507
rect 12149 44502 12150 44506
rect 11102 44442 12150 44502
rect 12400 44442 12401 44506
rect 12149 44441 12401 44442
rect 8878 44274 11168 44334
rect 8158 44215 8224 44250
rect 8113 44214 8481 44215
rect 8113 44142 8114 44214
rect 8480 44142 8481 44214
rect 10831 44154 10899 44155
rect 8113 44141 8481 44142
rect 9800 44026 10100 44154
rect 5950 43966 10100 44026
rect 10831 43976 10832 44154
rect 10898 43976 10899 44154
rect 11108 44053 11168 44274
rect 12574 44243 12634 45152
rect 13310 44633 13370 45152
rect 14046 44925 14106 45152
rect 13645 44906 14106 44925
rect 13645 44842 13683 44906
rect 13747 44842 13763 44906
rect 13827 44842 13843 44906
rect 13907 44842 13923 44906
rect 13987 44842 14003 44906
rect 14067 44888 14106 44906
rect 14067 44842 14105 44888
rect 13645 44823 14105 44842
rect 14782 44774 14842 45152
rect 14338 44758 14852 44774
rect 14338 44694 14361 44758
rect 14425 44694 14441 44758
rect 14505 44694 14521 44758
rect 14585 44694 14601 44758
rect 14665 44694 14681 44758
rect 14745 44694 14761 44758
rect 14825 44694 14852 44758
rect 14338 44682 14852 44694
rect 15518 44690 15578 45152
rect 16254 44856 16314 45152
rect 16619 44858 16685 44859
rect 16619 44856 16620 44858
rect 16254 44796 16620 44856
rect 16619 44794 16620 44796
rect 16684 44794 16685 44858
rect 16619 44793 16685 44794
rect 15873 44692 15939 44693
rect 15873 44690 15874 44692
rect 13035 44632 13475 44633
rect 13035 44568 13063 44632
rect 13127 44568 13143 44632
rect 13207 44568 13223 44632
rect 13287 44568 13303 44632
rect 13367 44568 13383 44632
rect 13447 44568 13475 44632
rect 15518 44630 15874 44690
rect 15873 44628 15874 44630
rect 15938 44628 15939 44692
rect 15873 44627 15939 44628
rect 13035 44567 13475 44568
rect 12843 44506 13141 44507
rect 12843 44438 12844 44506
rect 13140 44498 13141 44506
rect 13140 44438 16180 44498
rect 12843 44437 13141 44438
rect 12167 44242 12651 44243
rect 12167 44178 12177 44242
rect 12241 44178 12257 44242
rect 12321 44178 12337 44242
rect 12401 44178 12417 44242
rect 12481 44178 12497 44242
rect 12561 44178 12577 44242
rect 12641 44178 12651 44242
rect 12167 44177 12651 44178
rect 12574 44166 12634 44177
rect 10831 43975 10899 43976
rect 11001 44042 11229 44053
rect 9800 43873 10100 43966
rect 9799 43872 10107 43873
rect 4475 43828 4541 43829
rect 4475 43824 4476 43828
rect 3742 43764 4476 43824
rect 4540 43824 4541 43828
rect 4540 43764 4562 43824
rect 4475 43763 4541 43764
rect 9799 43624 9800 43872
rect 10106 43624 10107 43872
rect 9799 43623 10107 43624
rect 9800 42907 10100 43623
rect 9755 42906 10175 42907
rect 9755 42410 9756 42906
rect 10174 42410 10175 42906
rect 10838 42579 10898 43975
rect 11001 43738 11003 44042
rect 11227 43738 11229 44042
rect 11001 43727 11229 43738
rect 10838 42545 11123 42579
rect 10838 42412 10870 42545
rect 9755 42409 10175 42410
rect 1807 41838 2481 41839
rect 1807 41824 1808 41838
rect 200 41324 1808 41824
rect 200 34991 500 41324
rect 1807 41288 1808 41324
rect 2480 41824 2481 41838
rect 9800 41833 10100 42409
rect 10841 42401 10870 42412
rect 11094 42401 11123 42545
rect 10841 42367 11123 42401
rect 15775 42335 15841 42336
rect 15775 42271 15776 42335
rect 15840 42271 15841 42335
rect 15775 42270 15841 42271
rect 8529 41824 9031 41825
rect 2480 41719 8530 41824
rect 2480 41415 3865 41719
rect 5049 41415 8530 41719
rect 2480 41324 8530 41415
rect 9030 41324 9058 41824
rect 2480 41288 2481 41324
rect 8529 41323 9031 41324
rect 8700 41322 9000 41323
rect 9798 41313 10102 41833
rect 15059 41822 15679 41823
rect 15059 41336 15060 41822
rect 15678 41336 15679 41822
rect 15059 41335 15679 41336
rect 1807 41287 2481 41288
rect 9800 40419 10100 41313
rect 9800 40397 10515 40419
rect 9800 39933 10100 40397
rect 10507 39933 10515 40397
rect 9800 39911 10515 39933
rect 9800 37055 10100 39911
rect 15778 39072 15838 42270
rect 15959 42188 16025 42189
rect 15959 42124 15960 42188
rect 16024 42124 16025 42188
rect 15959 42123 16025 42124
rect 15962 39345 16022 42123
rect 16120 41248 16180 44438
rect 16990 42181 17050 45152
rect 17726 42352 17786 45152
rect 17712 42341 17808 42352
rect 17712 42277 17725 42341
rect 17789 42277 17808 42341
rect 17712 42264 17808 42277
rect 18462 42253 18522 45152
rect 19198 42375 19258 45152
rect 19934 44952 19994 45152
rect 20670 44952 20730 45152
rect 21406 42701 21466 45152
rect 22142 43893 22202 45152
rect 22878 44952 22938 45152
rect 21963 43870 22241 43893
rect 21963 43806 21990 43870
rect 22054 43806 22070 43870
rect 22134 43806 22150 43870
rect 22214 43806 22241 43870
rect 21963 43783 22241 43806
rect 21315 42699 21535 42701
rect 21315 42475 21353 42699
rect 21497 42475 21535 42699
rect 21315 42473 21535 42475
rect 19179 42348 19291 42375
rect 19179 42284 19203 42348
rect 19267 42284 19291 42348
rect 19179 42257 19291 42284
rect 18459 42233 18605 42253
rect 16987 42180 17053 42181
rect 16987 42116 16988 42180
rect 17052 42116 17053 42180
rect 16987 42115 17053 42116
rect 18459 42089 18460 42233
rect 18604 42089 18605 42233
rect 18459 42069 18605 42089
rect 16120 41226 17054 41248
rect 16120 41188 16952 41226
rect 16921 41162 16952 41188
rect 17016 41188 17054 41226
rect 17016 41162 17050 41188
rect 16921 41146 17050 41162
rect 16921 41082 16952 41146
rect 17016 41082 17050 41146
rect 16921 41066 17050 41082
rect 16921 41002 16952 41066
rect 17016 41002 17050 41066
rect 16921 40986 17050 41002
rect 16921 40922 16952 40986
rect 17016 40922 17050 40986
rect 23614 40941 23674 45152
rect 24350 44952 24410 45152
rect 23954 42385 24014 42388
rect 23935 42358 24047 42385
rect 23935 42294 23959 42358
rect 24023 42294 24047 42358
rect 23935 42267 24047 42294
rect 23936 42264 24042 42267
rect 16921 40906 17050 40922
rect 16921 40842 16952 40906
rect 17016 40842 17050 40906
rect 16921 40826 17050 40842
rect 16921 40762 16952 40826
rect 17016 40762 17050 40826
rect 16921 40745 17050 40762
rect 16990 40718 17050 40745
rect 23409 40905 23677 40941
rect 23409 40761 23431 40905
rect 23655 40761 23677 40905
rect 23409 40725 23677 40761
rect 23614 40718 23674 40725
rect 15955 39331 16033 39345
rect 15955 39267 15962 39331
rect 16026 39267 16033 39331
rect 15955 39253 16033 39267
rect 22151 39108 22327 39109
rect 18865 39074 19067 39103
rect 18865 39072 18894 39074
rect 15778 39012 18894 39072
rect 18836 38974 18894 39012
rect 18865 38930 18894 38974
rect 19038 38930 19067 39074
rect 18865 38901 19067 38930
rect 22151 38884 22167 39108
rect 22311 39010 22327 39108
rect 23982 39010 24042 42264
rect 24187 42146 24401 42167
rect 24187 42082 24222 42146
rect 24286 42082 24302 42146
rect 24366 42082 24401 42146
rect 24187 42061 24401 42082
rect 22311 38950 24048 39010
rect 22311 38884 22327 38950
rect 22151 38883 22327 38884
rect 15938 38813 16064 38836
rect 15938 38749 15962 38813
rect 16026 38749 16064 38813
rect 15938 38722 16064 38749
rect 15955 37281 16022 38722
rect 22137 37333 22323 37363
rect 18683 37298 18885 37327
rect 18683 37281 18712 37298
rect 15955 37209 18712 37281
rect 15955 37208 16015 37209
rect 18683 37154 18712 37209
rect 18856 37154 18885 37298
rect 22137 37189 22158 37333
rect 22302 37292 22323 37333
rect 24300 37292 24360 42061
rect 25086 38348 25146 45152
rect 25822 44952 25882 45152
rect 26558 44882 26618 45152
rect 25901 44833 26023 44857
rect 25901 44769 25930 44833
rect 25994 44769 26023 44833
rect 25901 44753 26023 44769
rect 25637 44657 25753 44693
rect 25901 44689 25930 44753
rect 25994 44689 26023 44753
rect 25901 44665 26023 44689
rect 26232 44822 26618 44882
rect 25637 44593 25663 44657
rect 25727 44593 25753 44657
rect 25637 44577 25753 44593
rect 25637 44513 25663 44577
rect 25727 44513 25753 44577
rect 25637 44477 25753 44513
rect 25692 43413 25752 44477
rect 25691 43408 25845 43413
rect 25691 43264 25696 43408
rect 25840 43264 25845 43408
rect 25691 43259 25845 43264
rect 25692 43250 25752 43259
rect 25962 41708 26022 44665
rect 26232 42277 26292 44822
rect 27294 44415 27354 45152
rect 27291 44414 27357 44415
rect 27291 44350 27292 44414
rect 27356 44350 27357 44414
rect 28030 44403 28090 45152
rect 27291 44349 27357 44350
rect 28005 44395 28127 44403
rect 28005 44331 28034 44395
rect 28098 44331 28127 44395
rect 28005 44315 28127 44331
rect 28005 44251 28034 44315
rect 28098 44251 28127 44315
rect 28005 44235 28127 44251
rect 28005 44171 28034 44235
rect 28098 44171 28127 44235
rect 28005 44155 28127 44171
rect 28005 44091 28034 44155
rect 28098 44091 28127 44155
rect 28005 44075 28127 44091
rect 28005 44011 28034 44075
rect 28098 44011 28127 44075
rect 28005 43995 28127 44011
rect 28005 43931 28034 43995
rect 28098 43931 28127 43995
rect 28005 43915 28127 43931
rect 28005 43851 28034 43915
rect 28098 43851 28127 43915
rect 28005 43843 28127 43851
rect 26199 42255 26343 42277
rect 26199 42191 26239 42255
rect 26303 42191 26343 42255
rect 26199 42175 26343 42191
rect 26199 42111 26239 42175
rect 26303 42111 26343 42175
rect 26199 42095 26343 42111
rect 26199 42031 26239 42095
rect 26303 42031 26343 42095
rect 26199 42015 26343 42031
rect 26199 41951 26239 42015
rect 26303 41951 26343 42015
rect 26199 41929 26343 41951
rect 26232 41924 26292 41929
rect 25962 41645 26028 41708
rect 25962 41633 26191 41645
rect 25962 41249 26008 41633
rect 26152 41249 26191 41633
rect 25962 41237 26191 41249
rect 25962 41228 26022 41237
rect 24604 38288 25146 38348
rect 22302 37232 24360 37292
rect 22302 37189 22323 37232
rect 22137 37159 22323 37189
rect 18683 37125 18885 37154
rect 9753 37054 10189 37055
rect 9753 36664 9754 37054
rect 10188 36664 10189 37054
rect 9753 36663 10189 36664
rect 9800 36321 10100 36663
rect 9800 36292 10489 36321
rect 9800 35428 10100 36292
rect 10481 35428 10489 36292
rect 9800 35399 10489 35428
rect 199 34986 1669 34991
rect 199 34122 222 34986
rect 1646 34122 1669 34986
rect 199 34117 1669 34122
rect 200 30699 500 34117
rect 200 30698 2363 30699
rect 200 29784 202 30698
rect 2362 29784 2363 30698
rect 200 29783 2363 29784
rect 200 6769 500 29783
rect 9800 26098 10100 35399
rect 24605 33933 24665 38288
rect 28766 35689 28826 45152
rect 29502 44950 29562 45152
rect 30238 44952 30298 45152
rect 30974 44952 31034 45152
rect 31710 44952 31770 45152
rect 29502 35717 29563 44950
rect 29489 35716 29595 35717
rect 28753 35688 28835 35689
rect 28753 35024 28754 35688
rect 28834 35024 28835 35688
rect 28753 35023 28835 35024
rect 29489 35014 29490 35716
rect 29594 35014 29595 35716
rect 29489 35013 29595 35014
rect 10863 33873 24665 33933
rect 10863 29867 10923 33873
rect 10355 29866 11159 29867
rect 10355 29428 10356 29866
rect 11158 29428 11159 29866
rect 10355 29427 11159 29428
rect 16281 26218 16711 26219
rect 16281 26098 16282 26218
rect 9800 25720 16282 26098
rect 200 6737 1017 6769
rect 200 6113 217 6737
rect 1001 6113 1017 6737
rect 200 6081 1017 6113
rect 200 1000 500 6081
rect 8165 1900 9399 1901
rect 8165 1554 8166 1900
rect 9398 1554 9399 1900
rect 8165 1553 9399 1554
rect 400 0 520 200
rect 4816 0 4936 200
rect 9232 0 9352 1553
rect 9800 1483 10100 25720
rect 16281 25712 16282 25720
rect 16710 25712 16711 26218
rect 16281 25711 16711 25712
rect 28747 6548 28847 6549
rect 28747 6074 28748 6548
rect 28846 6074 28847 6548
rect 29503 6545 29563 6546
rect 28747 6073 28847 6074
rect 29469 6544 29603 6545
rect 27367 4861 27643 4897
rect 27367 4808 27393 4861
rect 26934 4688 27393 4808
rect 25373 4027 25687 4049
rect 25373 3723 25378 4027
rect 25682 3723 25687 4027
rect 25373 3701 25687 3723
rect 19325 3593 19777 3631
rect 19325 3530 19359 3593
rect 18064 3449 19359 3530
rect 19743 3449 19777 3593
rect 18064 3411 19777 3449
rect 18064 3410 19754 3411
rect 13523 2792 13893 2793
rect 9800 1451 10589 1483
rect 9800 1067 10100 1451
rect 10583 1067 10589 1451
rect 9800 1035 10589 1067
rect 13523 1062 13524 2792
rect 13892 1062 13893 2792
rect 13523 1061 13893 1062
rect 9800 1000 10100 1035
rect 13648 0 13768 1061
rect 18064 0 18184 3410
rect 25452 888 25572 3701
rect 26934 1792 27054 4688
rect 27367 4637 27393 4688
rect 27617 4637 27643 4861
rect 27367 4601 27643 4637
rect 28766 2418 28826 6073
rect 29469 6062 29470 6544
rect 29602 6062 29603 6544
rect 29469 6061 29603 6062
rect 29503 3317 29563 6061
rect 29451 3312 29661 3317
rect 29451 3088 29484 3312
rect 29628 3088 29661 3312
rect 29451 3083 29661 3088
rect 29395 2432 29609 2457
rect 29395 2418 29430 2432
rect 28766 2358 29430 2418
rect 29395 2208 29430 2358
rect 29574 2208 29609 2432
rect 29395 2183 29609 2208
rect 31312 1792 31432 1800
rect 26934 1672 31440 1792
rect 26934 1660 27054 1672
rect 22480 768 25572 888
rect 26896 1050 30676 1078
rect 26896 986 30584 1050
rect 30648 986 30676 1050
rect 26896 958 30676 986
rect 22480 0 22600 768
rect 26896 0 27016 958
rect 31312 0 31432 1672
use cp  cp_0
timestamp 1712816020
transform 1 0 24094 0 1 7332
box 3292 -5232 7098 -1340
use Div  Div_0
timestamp 1712816020
transform 1 0 2194 0 -1 42140
box -670 -832 6794 -38
use divi_v1L  divi_v1L_0
timestamp 1713443771
transform 1 0 980 0 1 40194
box 974 -588 8440 630
use divider_tap  divider_tap_0
timestamp 1713443771
transform -1 0 23266 0 1 40038
box -402 448 6210 1246
use NFD_tap  NFD_tap_0
timestamp 1713443771
transform 0 -1 25184 1 0 36244
box 1330 -2334 7908 -1136
use Npfd  Npfd_0
timestamp 1713443771
transform -1 0 23222 0 1 38894
box 1024 -2182 4496 646
use Osc_v3_L  Osc_v3_L_0
timestamp 1712816020
transform -1 0 29132 0 1 3170
box 3508 -2212 9578 2934
use pfd_with_buffers_tap  pfd_with_buffers_tap_0
timestamp 1713443771
transform -1 0 17586 0 1 43836
box 1572 -1860 6566 514
use pll_integ  pll_integ_0 ~/pll/magic/pll_integ
timestamp 1713443771
transform 1 0 10796 0 1 27682
box -548 -20802 20064 5724
<< labels >>
flabel metal4 s 30974 44952 31034 45152 0 FreeSans 750 90 0 0 clk
port 1 nsew
flabel metal4 s 31710 44952 31770 45152 0 FreeSans 750 90 0 0 ena
port 2 nsew
flabel metal4 s 30238 44952 30298 45152 0 FreeSans 750 90 0 0 rst_n
port 3 nsew
flabel metal4 s 31312 0 31432 200 0 FreeSans 1500 0 0 0 ua[0]
port 4 nsew
flabel metal4 s 26896 0 27016 200 0 FreeSans 1500 0 0 0 ua[1]
port 5 nsew
flabel metal4 s 22480 0 22600 200 0 FreeSans 1500 0 0 0 ua[2]
port 6 nsew
flabel metal4 s 18064 0 18184 200 0 FreeSans 1500 0 0 0 ua[3]
port 7 nsew
flabel metal4 s 13648 0 13768 200 0 FreeSans 1500 0 0 0 ua[4]
port 8 nsew
flabel metal4 s 9232 0 9352 200 0 FreeSans 1500 0 0 0 ua[5]
port 9 nsew
flabel metal4 s 4816 0 4936 200 0 FreeSans 1500 0 0 0 ua[6]
port 10 nsew
flabel metal4 s 400 0 520 200 0 FreeSans 1500 0 0 0 ua[7]
port 11 nsew
flabel metal4 s 28766 44952 28826 45152 0 FreeSans 750 90 0 0 ui_in[1]
port 13 nsew
flabel metal4 s 28030 44952 28090 45152 0 FreeSans 750 90 0 0 ui_in[2]
port 14 nsew
flabel metal4 s 27294 44952 27354 45152 0 FreeSans 750 90 0 0 ui_in[3]
port 15 nsew
flabel metal4 s 26558 44952 26618 45152 0 FreeSans 750 90 0 0 ui_in[4]
port 16 nsew
flabel metal4 s 25822 44952 25882 45152 0 FreeSans 750 90 0 0 ui_in[5]
port 17 nsew
flabel metal4 s 25086 44952 25146 45152 0 FreeSans 750 90 0 0 ui_in[6]
port 18 nsew
flabel metal4 s 24350 44952 24410 45152 0 FreeSans 750 90 0 0 ui_in[7]
port 19 nsew
flabel metal4 s 23614 44952 23674 45152 0 FreeSans 750 90 0 0 uio_in[0]
port 20 nsew
flabel metal4 s 22878 44952 22938 45152 0 FreeSans 750 90 0 0 uio_in[1]
port 21 nsew
flabel metal4 s 22142 44952 22202 45152 0 FreeSans 750 90 0 0 uio_in[2]
port 22 nsew
flabel metal4 s 21406 44952 21466 45152 0 FreeSans 750 90 0 0 uio_in[3]
port 23 nsew
flabel metal4 s 20670 44952 20730 45152 0 FreeSans 750 90 0 0 uio_in[4]
port 24 nsew
flabel metal4 s 19934 44952 19994 45152 0 FreeSans 750 90 0 0 uio_in[5]
port 25 nsew
flabel metal4 s 19198 44952 19258 45152 0 FreeSans 750 90 0 0 uio_in[6]
port 26 nsew
flabel metal4 s 18462 44952 18522 45152 0 FreeSans 750 90 0 0 uio_in[7]
port 27 nsew
flabel metal4 s 5950 44952 6010 45152 0 FreeSans 750 90 0 0 uio_oe[0]
port 28 nsew
flabel metal4 s 5214 44952 5274 45152 0 FreeSans 750 90 0 0 uio_oe[1]
port 29 nsew
flabel metal4 s 4478 44952 4538 45152 0 FreeSans 750 90 0 0 uio_oe[2]
port 30 nsew
flabel metal4 s 3742 44952 3802 45152 0 FreeSans 750 90 0 0 uio_oe[3]
port 31 nsew
flabel metal4 s 3006 44952 3066 45152 0 FreeSans 750 90 0 0 uio_oe[4]
port 32 nsew
flabel metal4 s 2270 44952 2330 45152 0 FreeSans 750 90 0 0 uio_oe[5]
port 33 nsew
flabel metal4 s 1534 44952 1594 45152 0 FreeSans 750 90 0 0 uio_oe[6]
port 34 nsew
flabel metal4 s 798 44952 858 45152 0 FreeSans 750 90 0 0 uio_oe[7]
port 35 nsew
flabel metal4 s 11838 44952 11898 45152 0 FreeSans 750 90 0 0 uio_out[0]
port 36 nsew
flabel metal4 s 11102 44952 11162 45152 0 FreeSans 750 90 0 0 uio_out[1]
port 37 nsew
flabel metal4 s 10366 44952 10426 45152 0 FreeSans 750 90 0 0 uio_out[2]
port 38 nsew
flabel metal4 s 9630 44952 9690 45152 0 FreeSans 750 90 0 0 uio_out[3]
port 39 nsew
flabel metal4 s 8894 44952 8954 45152 0 FreeSans 750 90 0 0 uio_out[4]
port 40 nsew
flabel metal4 s 8158 44952 8218 45152 0 FreeSans 750 90 0 0 uio_out[5]
port 41 nsew
flabel metal4 s 7422 44952 7482 45152 0 FreeSans 750 90 0 0 uio_out[6]
port 42 nsew
flabel metal4 s 6686 44952 6746 45152 0 FreeSans 750 90 0 0 uio_out[7]
port 43 nsew
flabel metal4 s 17726 44952 17786 45152 0 FreeSans 750 90 0 0 uo_out[0]
port 44 nsew
flabel metal4 s 16990 44952 17050 45152 0 FreeSans 750 90 0 0 uo_out[1]
port 45 nsew
flabel metal4 s 16254 44952 16314 45152 0 FreeSans 750 90 0 0 uo_out[2]
port 46 nsew
flabel metal4 s 15518 44952 15578 45152 0 FreeSans 750 90 0 0 uo_out[3]
port 47 nsew
flabel metal4 s 14782 44952 14842 45152 0 FreeSans 750 90 0 0 uo_out[4]
port 48 nsew
flabel metal4 s 14046 44952 14106 45152 0 FreeSans 750 90 0 0 uo_out[5]
port 49 nsew
flabel metal4 s 13310 44952 13370 45152 0 FreeSans 750 90 0 0 uo_out[6]
port 50 nsew
flabel metal4 s 12574 44952 12634 45152 0 FreeSans 750 90 0 0 uo_out[7]
port 51 nsew
flabel metal4 s 200 1000 500 44152 1 FreeSans 2 0 0 0 VPWR
port 52 nsew
flabel metal4 9800 1000 10100 44152 1 FreeSans 2 0 0 0 VGND
port 53 n ground bidirectional
flabel metal4 s 29502 44952 29562 45152 0 FreeSans 750 90 0 0 ui_in[0]
port 12 nsew
<< properties >>
string FIXED_BBOX 0 0 32200 45152
<< end >>
