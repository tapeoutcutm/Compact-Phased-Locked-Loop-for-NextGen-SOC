magic
tech sky130A
magscale 1 2
timestamp 1713524523
<< nwell >>
rect 7674 -1760 7810 -1452
<< pwell >>
rect 1496 -1868 1642 -1866
rect 1496 -2026 1652 -1868
<< psubdiff >>
rect 1522 -1894 1616 -1892
rect 1522 -1929 1626 -1894
rect 1522 -1963 1557 -1929
rect 1591 -1963 1626 -1929
rect 1522 -2000 1626 -1963
<< nsubdiff >>
rect 7670 -1629 7774 -1570
rect 7670 -1663 7708 -1629
rect 7742 -1663 7774 -1629
rect 7670 -1718 7774 -1663
<< psubdiffcont >>
rect 1557 -1963 1591 -1929
<< nsubdiffcont >>
rect 7708 -1663 7742 -1629
<< locali >>
rect 7626 -1466 7772 -1458
rect 7626 -1472 7778 -1466
rect 7606 -1514 7778 -1472
rect 7672 -1629 7778 -1514
rect 7672 -1663 7708 -1629
rect 7742 -1663 7778 -1629
rect 7672 -1724 7778 -1663
rect 1402 -1765 1730 -1732
rect 1402 -1799 1415 -1765
rect 1449 -1799 1487 -1765
rect 1521 -1799 1730 -1765
rect 3450 -1772 3488 -1764
rect 1402 -1832 1730 -1799
rect 1936 -1794 1986 -1788
rect 1936 -1828 1944 -1794
rect 1978 -1828 1986 -1794
rect 3450 -1806 3452 -1772
rect 3486 -1778 3488 -1772
rect 5466 -1772 5504 -1764
rect 3486 -1806 3742 -1778
rect 3450 -1814 3742 -1806
rect 3958 -1788 4008 -1782
rect 3958 -1822 3966 -1788
rect 4000 -1822 4008 -1788
rect 5466 -1806 5468 -1772
rect 5502 -1780 5504 -1772
rect 7490 -1780 7528 -1772
rect 5502 -1806 5760 -1780
rect 5466 -1814 5760 -1806
rect 5982 -1788 6032 -1782
rect 3958 -1828 4008 -1822
rect 5982 -1822 5990 -1788
rect 6024 -1822 6032 -1788
rect 7490 -1814 7492 -1780
rect 7526 -1814 7528 -1780
rect 7490 -1822 7528 -1814
rect 5982 -1828 6032 -1822
rect 1936 -1834 1986 -1828
rect 1520 -1929 1624 -1894
rect 1520 -1963 1557 -1929
rect 1591 -1963 1624 -1929
rect 3044 -1906 3094 -1898
rect 3044 -1940 3052 -1906
rect 3086 -1940 3094 -1906
rect 3044 -1948 3094 -1940
rect 5066 -1906 5116 -1898
rect 5066 -1940 5074 -1906
rect 5108 -1940 5116 -1906
rect 5066 -1948 5116 -1940
rect 7090 -1906 7140 -1898
rect 7090 -1940 7098 -1906
rect 7132 -1940 7140 -1906
rect 7090 -1948 7140 -1940
rect 1520 -2018 1624 -1963
rect 1520 -2056 1686 -2018
<< viali >>
rect 1415 -1799 1449 -1765
rect 1487 -1799 1521 -1765
rect 1944 -1828 1978 -1794
rect 3452 -1806 3486 -1772
rect 3966 -1822 4000 -1788
rect 5468 -1806 5502 -1772
rect 5990 -1822 6024 -1788
rect 7492 -1814 7526 -1780
rect 3052 -1940 3086 -1906
rect 5074 -1940 5108 -1906
rect 7098 -1940 7132 -1906
<< metal1 >>
rect 1330 -1440 1530 -1136
rect 2960 -1319 3160 -1162
rect 2960 -1362 3000 -1319
rect 2982 -1371 3000 -1362
rect 3052 -1371 3064 -1319
rect 3116 -1362 3160 -1319
rect 4982 -1327 5182 -1168
rect 3116 -1371 3134 -1362
rect 4982 -1368 5030 -1327
rect 2982 -1386 3134 -1371
rect 5012 -1379 5030 -1368
rect 5082 -1379 5094 -1327
rect 5146 -1368 5182 -1327
rect 7000 -1333 7200 -1166
rect 7000 -1366 7046 -1333
rect 5146 -1379 5164 -1368
rect 5012 -1394 5164 -1379
rect 7028 -1385 7046 -1366
rect 7098 -1385 7110 -1333
rect 7162 -1366 7200 -1333
rect 7162 -1385 7180 -1366
rect 7028 -1400 7180 -1385
rect 1330 -1534 1740 -1440
rect 5022 -1581 5148 -1576
rect 3000 -1595 3126 -1590
rect 3000 -1647 3037 -1595
rect 3089 -1647 3126 -1595
rect 5022 -1633 5059 -1581
rect 5111 -1633 5148 -1581
rect 5022 -1638 5148 -1633
rect 7044 -1587 7170 -1582
rect 3000 -1652 3126 -1647
rect 1334 -1726 1534 -1686
rect 1334 -1765 1546 -1726
rect 1334 -1799 1415 -1765
rect 1449 -1799 1487 -1765
rect 1521 -1799 1546 -1765
rect 1974 -1782 2928 -1780
rect 1334 -1838 1546 -1799
rect 1924 -1786 2928 -1782
rect 1924 -1794 2853 -1786
rect 1924 -1828 1944 -1794
rect 1978 -1828 2853 -1794
rect 1924 -1838 2853 -1828
rect 2905 -1838 2928 -1786
rect 1334 -1886 1534 -1838
rect 1924 -1840 2928 -1838
rect 1974 -1842 2928 -1840
rect 2830 -1844 2928 -1842
rect 3026 -1902 3106 -1652
rect 3444 -1754 3494 -1752
rect 3374 -1764 3494 -1754
rect 3374 -1816 3386 -1764
rect 3438 -1772 3494 -1764
rect 3438 -1806 3452 -1772
rect 3486 -1806 3494 -1772
rect 4860 -1766 4958 -1760
rect 3438 -1816 3494 -1806
rect 3374 -1826 3494 -1816
rect 3946 -1786 4020 -1776
rect 4860 -1786 4883 -1766
rect 3946 -1788 4883 -1786
rect 3946 -1822 3966 -1788
rect 4000 -1818 4883 -1788
rect 4935 -1818 4958 -1766
rect 4000 -1822 4958 -1818
rect 3946 -1824 4958 -1822
rect 3946 -1832 4876 -1824
rect 3946 -1834 4020 -1832
rect 3032 -1906 3106 -1902
rect 3032 -1940 3052 -1906
rect 3086 -1940 3106 -1906
rect 3032 -1954 3106 -1940
rect 5054 -1892 5120 -1638
rect 7044 -1639 7081 -1587
rect 7133 -1639 7170 -1587
rect 7044 -1644 7170 -1639
rect 5396 -1762 5510 -1752
rect 5396 -1814 5408 -1762
rect 5460 -1772 5510 -1762
rect 5460 -1806 5468 -1772
rect 5502 -1806 5510 -1772
rect 5460 -1814 5510 -1806
rect 5396 -1824 5510 -1814
rect 5460 -1826 5510 -1824
rect 5970 -1782 6044 -1776
rect 6924 -1778 7022 -1772
rect 6924 -1782 6947 -1778
rect 5970 -1788 6947 -1782
rect 5970 -1822 5990 -1788
rect 6024 -1822 6947 -1788
rect 5970 -1830 6947 -1822
rect 6999 -1830 7022 -1778
rect 5970 -1832 7022 -1830
rect 5970 -1834 6044 -1832
rect 6924 -1836 7022 -1832
rect 5054 -1906 5128 -1892
rect 7076 -1906 7152 -1644
rect 7428 -1770 7534 -1760
rect 7428 -1822 7440 -1770
rect 7492 -1780 7534 -1770
rect 7526 -1814 7534 -1780
rect 7492 -1822 7534 -1814
rect 7428 -1832 7534 -1822
rect 7484 -1834 7534 -1832
rect 5054 -1940 5074 -1906
rect 5108 -1940 5128 -1906
rect 5054 -1954 5128 -1940
rect 7078 -1940 7098 -1906
rect 7132 -1940 7152 -1906
rect 7078 -1954 7152 -1940
rect 7550 -2006 7636 -1998
rect 7550 -2080 7904 -2006
rect 7708 -2134 7904 -2080
rect 7708 -2334 7908 -2134
<< via1 >>
rect 3000 -1371 3052 -1319
rect 3064 -1371 3116 -1319
rect 5030 -1379 5082 -1327
rect 5094 -1379 5146 -1327
rect 7046 -1385 7098 -1333
rect 7110 -1385 7162 -1333
rect 3037 -1647 3089 -1595
rect 5059 -1633 5111 -1581
rect 2853 -1838 2905 -1786
rect 3386 -1816 3438 -1764
rect 4883 -1818 4935 -1766
rect 7081 -1639 7133 -1587
rect 5408 -1814 5460 -1762
rect 6947 -1830 6999 -1778
rect 7440 -1822 7492 -1770
<< metal2 >>
rect 2992 -1319 3124 -1294
rect 2992 -1371 3000 -1319
rect 3052 -1371 3064 -1319
rect 3116 -1371 3124 -1319
rect 2992 -1378 3124 -1371
rect 5022 -1327 5154 -1302
rect 2992 -1396 3126 -1378
rect 2996 -1594 3126 -1396
rect 5022 -1379 5030 -1327
rect 5082 -1379 5094 -1327
rect 5146 -1379 5154 -1327
rect 5022 -1404 5154 -1379
rect 7038 -1333 7170 -1308
rect 7038 -1385 7046 -1333
rect 7098 -1385 7110 -1333
rect 7162 -1385 7170 -1333
rect 5038 -1566 5132 -1404
rect 7038 -1410 7170 -1385
rect 5032 -1581 5138 -1566
rect 3010 -1595 3116 -1594
rect 3010 -1647 3037 -1595
rect 3089 -1647 3116 -1595
rect 3010 -1662 3116 -1647
rect 5032 -1633 5059 -1581
rect 5111 -1633 5138 -1581
rect 7050 -1584 7162 -1410
rect 5032 -1648 5138 -1633
rect 7054 -1587 7160 -1584
rect 7054 -1639 7081 -1587
rect 7133 -1639 7160 -1587
rect 7054 -1654 7160 -1639
rect 3384 -1756 3440 -1744
rect 3024 -1768 3106 -1756
rect 3372 -1764 3440 -1756
rect 3372 -1768 3386 -1764
rect 2910 -1770 3386 -1768
rect 2840 -1786 3386 -1770
rect 2840 -1838 2853 -1786
rect 2905 -1816 3386 -1786
rect 3438 -1816 3440 -1764
rect 2905 -1834 3440 -1816
rect 4870 -1760 4948 -1750
rect 5406 -1760 5462 -1742
rect 4870 -1762 5462 -1760
rect 4870 -1766 5408 -1762
rect 4870 -1818 4883 -1766
rect 4935 -1814 5408 -1766
rect 5460 -1814 5462 -1762
rect 4935 -1818 5462 -1814
rect 4870 -1834 4948 -1818
rect 5406 -1834 5462 -1818
rect 6934 -1768 7012 -1762
rect 6934 -1770 7356 -1768
rect 7438 -1770 7494 -1750
rect 6934 -1778 7440 -1770
rect 6934 -1830 6947 -1778
rect 6999 -1822 7440 -1778
rect 7492 -1822 7494 -1770
rect 6999 -1830 7494 -1822
rect 6934 -1832 7494 -1830
rect 6934 -1834 7356 -1832
rect 2905 -1838 2928 -1834
rect 2840 -1844 2928 -1838
rect 3026 -1836 3440 -1834
rect 3026 -1844 3106 -1836
rect 2840 -1854 2918 -1844
rect 6934 -1846 7012 -1834
rect 7438 -1842 7494 -1832
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1712078602
transform 1 0 3588 0 1 -2034
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_1
timestamp 1712078602
transform 1 0 5612 0 1 -2034
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_2  x1 ~/pll/magic/divider
timestamp 1713423503
transform 1 0 1658 0 1 -2034
box -38 -48 1970 592
use sky130_fd_sc_hd__dfxbp_2  x2
timestamp 1713423503
transform 1 0 3680 0 1 -2034
box -38 -48 1970 592
use sky130_fd_sc_hd__dfxbp_2  x3
timestamp 1713423503
transform 1 0 5704 0 1 -2034
box -38 -48 1970 592
<< labels >>
flabel metal1 s 7708 -2334 7908 -2134 0 FreeSans 500 0 0 0 VSS
port 1 nsew
flabel metal1 s 7000 -1366 7200 -1166 0 FreeSans 500 0 0 0 f0_8
port 2 nsew
flabel metal1 s 4982 -1368 5182 -1168 0 FreeSans 500 0 0 0 f0_4
port 3 nsew
flabel metal1 s 2960 -1362 3160 -1162 0 FreeSans 500 0 0 0 f0_2
port 4 nsew
flabel metal1 s 1330 -1336 1530 -1136 0 FreeSans 500 0 0 0 VDD
port 5 nsew
flabel metal1 s 1334 -1886 1534 -1686 0 FreeSans 500 0 0 0 clk
port 6 nsew
<< end >>
