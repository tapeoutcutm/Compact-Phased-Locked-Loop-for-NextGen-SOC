magic
tech sky130A
magscale 1 2
timestamp 1712816020
<< nwell >>
rect -479 -419 479 419
<< pmos >>
rect -283 -200 -133 200
rect -75 -200 75 200
rect 133 -200 283 200
<< pdiff >>
rect -341 187 -283 200
rect -341 153 -329 187
rect -295 153 -283 187
rect -341 119 -283 153
rect -341 85 -329 119
rect -295 85 -283 119
rect -341 51 -283 85
rect -341 17 -329 51
rect -295 17 -283 51
rect -341 -17 -283 17
rect -341 -51 -329 -17
rect -295 -51 -283 -17
rect -341 -85 -283 -51
rect -341 -119 -329 -85
rect -295 -119 -283 -85
rect -341 -153 -283 -119
rect -341 -187 -329 -153
rect -295 -187 -283 -153
rect -341 -200 -283 -187
rect -133 187 -75 200
rect -133 153 -121 187
rect -87 153 -75 187
rect -133 119 -75 153
rect -133 85 -121 119
rect -87 85 -75 119
rect -133 51 -75 85
rect -133 17 -121 51
rect -87 17 -75 51
rect -133 -17 -75 17
rect -133 -51 -121 -17
rect -87 -51 -75 -17
rect -133 -85 -75 -51
rect -133 -119 -121 -85
rect -87 -119 -75 -85
rect -133 -153 -75 -119
rect -133 -187 -121 -153
rect -87 -187 -75 -153
rect -133 -200 -75 -187
rect 75 187 133 200
rect 75 153 87 187
rect 121 153 133 187
rect 75 119 133 153
rect 75 85 87 119
rect 121 85 133 119
rect 75 51 133 85
rect 75 17 87 51
rect 121 17 133 51
rect 75 -17 133 17
rect 75 -51 87 -17
rect 121 -51 133 -17
rect 75 -85 133 -51
rect 75 -119 87 -85
rect 121 -119 133 -85
rect 75 -153 133 -119
rect 75 -187 87 -153
rect 121 -187 133 -153
rect 75 -200 133 -187
rect 283 187 341 200
rect 283 153 295 187
rect 329 153 341 187
rect 283 119 341 153
rect 283 85 295 119
rect 329 85 341 119
rect 283 51 341 85
rect 283 17 295 51
rect 329 17 341 51
rect 283 -17 341 17
rect 283 -51 295 -17
rect 329 -51 341 -17
rect 283 -85 341 -51
rect 283 -119 295 -85
rect 329 -119 341 -85
rect 283 -153 341 -119
rect 283 -187 295 -153
rect 329 -187 341 -153
rect 283 -200 341 -187
<< pdiffc >>
rect -329 153 -295 187
rect -329 85 -295 119
rect -329 17 -295 51
rect -329 -51 -295 -17
rect -329 -119 -295 -85
rect -329 -187 -295 -153
rect -121 153 -87 187
rect -121 85 -87 119
rect -121 17 -87 51
rect -121 -51 -87 -17
rect -121 -119 -87 -85
rect -121 -187 -87 -153
rect 87 153 121 187
rect 87 85 121 119
rect 87 17 121 51
rect 87 -51 121 -17
rect 87 -119 121 -85
rect 87 -187 121 -153
rect 295 153 329 187
rect 295 85 329 119
rect 295 17 329 51
rect 295 -51 329 -17
rect 295 -119 329 -85
rect 295 -187 329 -153
<< nsubdiff >>
rect -443 349 -323 383
rect -289 349 -255 383
rect -221 349 -187 383
rect -153 349 -119 383
rect -85 349 -51 383
rect -17 349 17 383
rect 51 349 85 383
rect 119 349 153 383
rect 187 349 221 383
rect 255 349 289 383
rect 323 349 443 383
rect -443 255 -409 349
rect -443 187 -409 221
rect 409 255 443 349
rect -443 119 -409 153
rect -443 51 -409 85
rect -443 -17 -409 17
rect -443 -85 -409 -51
rect -443 -153 -409 -119
rect -443 -221 -409 -187
rect 409 187 443 221
rect 409 119 443 153
rect 409 51 443 85
rect 409 -17 443 17
rect 409 -85 443 -51
rect 409 -153 443 -119
rect -443 -349 -409 -255
rect 409 -221 443 -187
rect 409 -349 443 -255
rect -443 -383 -323 -349
rect -289 -383 -255 -349
rect -221 -383 -187 -349
rect -153 -383 -119 -349
rect -85 -383 -51 -349
rect -17 -383 17 -349
rect 51 -383 85 -349
rect 119 -383 153 -349
rect 187 -383 221 -349
rect 255 -383 289 -349
rect 323 -383 443 -349
<< nsubdiffcont >>
rect -323 349 -289 383
rect -255 349 -221 383
rect -187 349 -153 383
rect -119 349 -85 383
rect -51 349 -17 383
rect 17 349 51 383
rect 85 349 119 383
rect 153 349 187 383
rect 221 349 255 383
rect 289 349 323 383
rect -443 221 -409 255
rect 409 221 443 255
rect -443 153 -409 187
rect -443 85 -409 119
rect -443 17 -409 51
rect -443 -51 -409 -17
rect -443 -119 -409 -85
rect -443 -187 -409 -153
rect 409 153 443 187
rect 409 85 443 119
rect 409 17 443 51
rect 409 -51 443 -17
rect 409 -119 443 -85
rect 409 -187 443 -153
rect -443 -255 -409 -221
rect 409 -255 443 -221
rect -323 -383 -289 -349
rect -255 -383 -221 -349
rect -187 -383 -153 -349
rect -119 -383 -85 -349
rect -51 -383 -17 -349
rect 17 -383 51 -349
rect 85 -383 119 -349
rect 153 -383 187 -349
rect 221 -383 255 -349
rect 289 -383 323 -349
<< poly >>
rect -283 281 -133 297
rect -283 247 -259 281
rect -225 247 -191 281
rect -157 247 -133 281
rect -283 200 -133 247
rect -75 281 75 297
rect -75 247 -51 281
rect -17 247 17 281
rect 51 247 75 281
rect -75 200 75 247
rect 133 281 283 297
rect 133 247 157 281
rect 191 247 225 281
rect 259 247 283 281
rect 133 200 283 247
rect -283 -247 -133 -200
rect -283 -281 -259 -247
rect -225 -281 -191 -247
rect -157 -281 -133 -247
rect -283 -297 -133 -281
rect -75 -247 75 -200
rect -75 -281 -51 -247
rect -17 -281 17 -247
rect 51 -281 75 -247
rect -75 -297 75 -281
rect 133 -247 283 -200
rect 133 -281 157 -247
rect 191 -281 225 -247
rect 259 -281 283 -247
rect 133 -297 283 -281
<< polycont >>
rect -259 247 -225 281
rect -191 247 -157 281
rect -51 247 -17 281
rect 17 247 51 281
rect 157 247 191 281
rect 225 247 259 281
rect -259 -281 -225 -247
rect -191 -281 -157 -247
rect -51 -281 -17 -247
rect 17 -281 51 -247
rect 157 -281 191 -247
rect 225 -281 259 -247
<< locali >>
rect -443 349 -323 383
rect -289 349 -255 383
rect -221 349 -187 383
rect -153 349 -119 383
rect -85 349 -51 383
rect -17 349 17 383
rect 51 349 85 383
rect 119 349 153 383
rect 187 349 221 383
rect 255 349 289 383
rect 323 349 443 383
rect -443 255 -409 349
rect -283 247 -261 281
rect -225 247 -191 281
rect -155 247 -133 281
rect -75 247 -53 281
rect -17 247 17 281
rect 53 247 75 281
rect 133 247 155 281
rect 191 247 225 281
rect 261 247 283 281
rect 409 255 443 349
rect -443 187 -409 221
rect -443 119 -409 153
rect -443 51 -409 85
rect -443 -17 -409 17
rect -443 -85 -409 -51
rect -443 -153 -409 -119
rect -443 -221 -409 -187
rect -329 187 -295 204
rect -329 119 -295 127
rect -329 51 -295 55
rect -329 -55 -295 -51
rect -329 -127 -295 -119
rect -329 -204 -295 -187
rect -121 187 -87 204
rect -121 119 -87 127
rect -121 51 -87 55
rect -121 -55 -87 -51
rect -121 -127 -87 -119
rect -121 -204 -87 -187
rect 87 187 121 204
rect 87 119 121 127
rect 87 51 121 55
rect 87 -55 121 -51
rect 87 -127 121 -119
rect 87 -204 121 -187
rect 295 187 329 204
rect 295 119 329 127
rect 295 51 329 55
rect 295 -55 329 -51
rect 295 -127 329 -119
rect 295 -204 329 -187
rect 409 187 443 221
rect 409 119 443 153
rect 409 51 443 85
rect 409 -17 443 17
rect 409 -85 443 -51
rect 409 -153 443 -119
rect 409 -221 443 -187
rect -443 -349 -409 -255
rect -283 -281 -261 -247
rect -225 -281 -191 -247
rect -155 -281 -133 -247
rect -75 -281 -53 -247
rect -17 -281 17 -247
rect 53 -281 75 -247
rect 133 -281 155 -247
rect 191 -281 225 -247
rect 261 -281 283 -247
rect 409 -349 443 -255
rect -443 -383 -323 -349
rect -289 -383 -255 -349
rect -221 -383 -187 -349
rect -153 -383 -119 -349
rect -85 -383 -51 -349
rect -17 -383 17 -349
rect 51 -383 85 -349
rect 119 -383 153 -349
rect 187 -383 221 -349
rect 255 -383 289 -349
rect 323 -383 443 -349
<< viali >>
rect -261 247 -259 281
rect -259 247 -227 281
rect -189 247 -157 281
rect -157 247 -155 281
rect -53 247 -51 281
rect -51 247 -19 281
rect 19 247 51 281
rect 51 247 53 281
rect 155 247 157 281
rect 157 247 189 281
rect 227 247 259 281
rect 259 247 261 281
rect -329 153 -295 161
rect -329 127 -295 153
rect -329 85 -295 89
rect -329 55 -295 85
rect -329 -17 -295 17
rect -329 -85 -295 -55
rect -329 -89 -295 -85
rect -329 -153 -295 -127
rect -329 -161 -295 -153
rect -121 153 -87 161
rect -121 127 -87 153
rect -121 85 -87 89
rect -121 55 -87 85
rect -121 -17 -87 17
rect -121 -85 -87 -55
rect -121 -89 -87 -85
rect -121 -153 -87 -127
rect -121 -161 -87 -153
rect 87 153 121 161
rect 87 127 121 153
rect 87 85 121 89
rect 87 55 121 85
rect 87 -17 121 17
rect 87 -85 121 -55
rect 87 -89 121 -85
rect 87 -153 121 -127
rect 87 -161 121 -153
rect 295 153 329 161
rect 295 127 329 153
rect 295 85 329 89
rect 295 55 329 85
rect 295 -17 329 17
rect 295 -85 329 -55
rect 295 -89 329 -85
rect 295 -153 329 -127
rect 295 -161 329 -153
rect -261 -281 -259 -247
rect -259 -281 -227 -247
rect -189 -281 -157 -247
rect -157 -281 -155 -247
rect -53 -281 -51 -247
rect -51 -281 -19 -247
rect 19 -281 51 -247
rect 51 -281 53 -247
rect 155 -281 157 -247
rect 157 -281 189 -247
rect 227 -281 259 -247
rect 259 -281 261 -247
<< metal1 >>
rect -279 281 -137 287
rect -279 247 -261 281
rect -227 247 -189 281
rect -155 247 -137 281
rect -279 241 -137 247
rect -71 281 71 287
rect -71 247 -53 281
rect -19 247 19 281
rect 53 247 71 281
rect -71 241 71 247
rect 137 281 279 287
rect 137 247 155 281
rect 189 247 227 281
rect 261 247 279 281
rect 137 241 279 247
rect -335 161 -289 200
rect -335 127 -329 161
rect -295 127 -289 161
rect -335 89 -289 127
rect -335 55 -329 89
rect -295 55 -289 89
rect -335 17 -289 55
rect -335 -17 -329 17
rect -295 -17 -289 17
rect -335 -55 -289 -17
rect -335 -89 -329 -55
rect -295 -89 -289 -55
rect -335 -127 -289 -89
rect -335 -161 -329 -127
rect -295 -161 -289 -127
rect -335 -200 -289 -161
rect -127 161 -81 200
rect -127 127 -121 161
rect -87 127 -81 161
rect -127 89 -81 127
rect -127 55 -121 89
rect -87 55 -81 89
rect -127 17 -81 55
rect -127 -17 -121 17
rect -87 -17 -81 17
rect -127 -55 -81 -17
rect -127 -89 -121 -55
rect -87 -89 -81 -55
rect -127 -127 -81 -89
rect -127 -161 -121 -127
rect -87 -161 -81 -127
rect -127 -200 -81 -161
rect 81 161 127 200
rect 81 127 87 161
rect 121 127 127 161
rect 81 89 127 127
rect 81 55 87 89
rect 121 55 127 89
rect 81 17 127 55
rect 81 -17 87 17
rect 121 -17 127 17
rect 81 -55 127 -17
rect 81 -89 87 -55
rect 121 -89 127 -55
rect 81 -127 127 -89
rect 81 -161 87 -127
rect 121 -161 127 -127
rect 81 -200 127 -161
rect 289 161 335 200
rect 289 127 295 161
rect 329 127 335 161
rect 289 89 335 127
rect 289 55 295 89
rect 329 55 335 89
rect 289 17 335 55
rect 289 -17 295 17
rect 329 -17 335 17
rect 289 -55 335 -17
rect 289 -89 295 -55
rect 329 -89 335 -55
rect 289 -127 335 -89
rect 289 -161 295 -127
rect 329 -161 335 -127
rect 289 -200 335 -161
rect -279 -247 -137 -241
rect -279 -281 -261 -247
rect -227 -281 -189 -247
rect -155 -281 -137 -247
rect -279 -287 -137 -281
rect -71 -247 71 -241
rect -71 -281 -53 -247
rect -19 -281 19 -247
rect 53 -281 71 -247
rect -71 -287 71 -281
rect 137 -247 279 -241
rect 137 -281 155 -247
rect 189 -281 227 -247
rect 261 -281 279 -247
rect 137 -287 279 -281
<< properties >>
string FIXED_BBOX -426 -366 426 366
<< end >>
