magic
tech sky130A
magscale 1 2
timestamp 1712737205
<< pwell >>
rect -375 -525 375 525
<< nmos >>
rect -189 -325 -29 325
rect 29 -325 189 325
<< ndiff >>
rect -247 289 -189 325
rect -247 255 -235 289
rect -201 255 -189 289
rect -247 221 -189 255
rect -247 187 -235 221
rect -201 187 -189 221
rect -247 153 -189 187
rect -247 119 -235 153
rect -201 119 -189 153
rect -247 85 -189 119
rect -247 51 -235 85
rect -201 51 -189 85
rect -247 17 -189 51
rect -247 -17 -235 17
rect -201 -17 -189 17
rect -247 -51 -189 -17
rect -247 -85 -235 -51
rect -201 -85 -189 -51
rect -247 -119 -189 -85
rect -247 -153 -235 -119
rect -201 -153 -189 -119
rect -247 -187 -189 -153
rect -247 -221 -235 -187
rect -201 -221 -189 -187
rect -247 -255 -189 -221
rect -247 -289 -235 -255
rect -201 -289 -189 -255
rect -247 -325 -189 -289
rect -29 289 29 325
rect -29 255 -17 289
rect 17 255 29 289
rect -29 221 29 255
rect -29 187 -17 221
rect 17 187 29 221
rect -29 153 29 187
rect -29 119 -17 153
rect 17 119 29 153
rect -29 85 29 119
rect -29 51 -17 85
rect 17 51 29 85
rect -29 17 29 51
rect -29 -17 -17 17
rect 17 -17 29 17
rect -29 -51 29 -17
rect -29 -85 -17 -51
rect 17 -85 29 -51
rect -29 -119 29 -85
rect -29 -153 -17 -119
rect 17 -153 29 -119
rect -29 -187 29 -153
rect -29 -221 -17 -187
rect 17 -221 29 -187
rect -29 -255 29 -221
rect -29 -289 -17 -255
rect 17 -289 29 -255
rect -29 -325 29 -289
rect 189 289 247 325
rect 189 255 201 289
rect 235 255 247 289
rect 189 221 247 255
rect 189 187 201 221
rect 235 187 247 221
rect 189 153 247 187
rect 189 119 201 153
rect 235 119 247 153
rect 189 85 247 119
rect 189 51 201 85
rect 235 51 247 85
rect 189 17 247 51
rect 189 -17 201 17
rect 235 -17 247 17
rect 189 -51 247 -17
rect 189 -85 201 -51
rect 235 -85 247 -51
rect 189 -119 247 -85
rect 189 -153 201 -119
rect 235 -153 247 -119
rect 189 -187 247 -153
rect 189 -221 201 -187
rect 235 -221 247 -187
rect 189 -255 247 -221
rect 189 -289 201 -255
rect 235 -289 247 -255
rect 189 -325 247 -289
<< ndiffc >>
rect -235 255 -201 289
rect -235 187 -201 221
rect -235 119 -201 153
rect -235 51 -201 85
rect -235 -17 -201 17
rect -235 -85 -201 -51
rect -235 -153 -201 -119
rect -235 -221 -201 -187
rect -235 -289 -201 -255
rect -17 255 17 289
rect -17 187 17 221
rect -17 119 17 153
rect -17 51 17 85
rect -17 -17 17 17
rect -17 -85 17 -51
rect -17 -153 17 -119
rect -17 -221 17 -187
rect -17 -289 17 -255
rect 201 255 235 289
rect 201 187 235 221
rect 201 119 235 153
rect 201 51 235 85
rect 201 -17 235 17
rect 201 -85 235 -51
rect 201 -153 235 -119
rect 201 -221 235 -187
rect 201 -289 235 -255
<< psubdiff >>
rect -349 465 -221 499
rect -187 465 -153 499
rect -119 465 -85 499
rect -51 465 -17 499
rect 17 465 51 499
rect 85 465 119 499
rect 153 465 187 499
rect 221 465 349 499
rect -349 391 -315 465
rect -349 323 -315 357
rect 315 391 349 465
rect -349 255 -315 289
rect -349 187 -315 221
rect -349 119 -315 153
rect -349 51 -315 85
rect -349 -17 -315 17
rect -349 -85 -315 -51
rect -349 -153 -315 -119
rect -349 -221 -315 -187
rect -349 -289 -315 -255
rect -349 -357 -315 -323
rect 315 323 349 357
rect 315 255 349 289
rect 315 187 349 221
rect 315 119 349 153
rect 315 51 349 85
rect 315 -17 349 17
rect 315 -85 349 -51
rect 315 -153 349 -119
rect 315 -221 349 -187
rect 315 -289 349 -255
rect -349 -465 -315 -391
rect 315 -357 349 -323
rect 315 -465 349 -391
rect -349 -499 -221 -465
rect -187 -499 -153 -465
rect -119 -499 -85 -465
rect -51 -499 -17 -465
rect 17 -499 51 -465
rect 85 -499 119 -465
rect 153 -499 187 -465
rect 221 -499 349 -465
<< psubdiffcont >>
rect -221 465 -187 499
rect -153 465 -119 499
rect -85 465 -51 499
rect -17 465 17 499
rect 51 465 85 499
rect 119 465 153 499
rect 187 465 221 499
rect -349 357 -315 391
rect 315 357 349 391
rect -349 289 -315 323
rect -349 221 -315 255
rect -349 153 -315 187
rect -349 85 -315 119
rect -349 17 -315 51
rect -349 -51 -315 -17
rect -349 -119 -315 -85
rect -349 -187 -315 -153
rect -349 -255 -315 -221
rect -349 -323 -315 -289
rect 315 289 349 323
rect 315 221 349 255
rect 315 153 349 187
rect 315 85 349 119
rect 315 17 349 51
rect 315 -51 349 -17
rect 315 -119 349 -85
rect 315 -187 349 -153
rect 315 -255 349 -221
rect 315 -323 349 -289
rect -349 -391 -315 -357
rect 315 -391 349 -357
rect -221 -499 -187 -465
rect -153 -499 -119 -465
rect -85 -499 -51 -465
rect -17 -499 17 -465
rect 51 -499 85 -465
rect 119 -499 153 -465
rect 187 -499 221 -465
<< poly >>
rect -189 397 -29 413
rect -189 363 -160 397
rect -126 363 -92 397
rect -58 363 -29 397
rect -189 325 -29 363
rect 29 397 189 413
rect 29 363 58 397
rect 92 363 126 397
rect 160 363 189 397
rect 29 325 189 363
rect -189 -363 -29 -325
rect -189 -397 -160 -363
rect -126 -397 -92 -363
rect -58 -397 -29 -363
rect -189 -413 -29 -397
rect 29 -363 189 -325
rect 29 -397 58 -363
rect 92 -397 126 -363
rect 160 -397 189 -363
rect 29 -413 189 -397
<< polycont >>
rect -160 363 -126 397
rect -92 363 -58 397
rect 58 363 92 397
rect 126 363 160 397
rect -160 -397 -126 -363
rect -92 -397 -58 -363
rect 58 -397 92 -363
rect 126 -397 160 -363
<< locali >>
rect -349 465 -221 499
rect -187 465 -153 499
rect -119 465 -85 499
rect -51 465 -17 499
rect 17 465 51 499
rect 85 465 119 499
rect 153 465 187 499
rect 221 465 349 499
rect -349 391 -315 465
rect -189 363 -162 397
rect -126 363 -92 397
rect -56 363 -29 397
rect 29 363 56 397
rect 92 363 126 397
rect 162 363 189 397
rect 315 391 349 465
rect -349 323 -315 357
rect -349 255 -315 289
rect -349 187 -315 221
rect -349 119 -315 153
rect -349 51 -315 85
rect -349 -17 -315 17
rect -349 -85 -315 -51
rect -349 -153 -315 -119
rect -349 -221 -315 -187
rect -349 -289 -315 -255
rect -349 -357 -315 -323
rect -235 305 -201 329
rect -235 233 -201 255
rect -235 161 -201 187
rect -235 89 -201 119
rect -235 17 -201 51
rect -235 -51 -201 -17
rect -235 -119 -201 -89
rect -235 -187 -201 -161
rect -235 -255 -201 -233
rect -235 -329 -201 -305
rect -17 305 17 329
rect -17 233 17 255
rect -17 161 17 187
rect -17 89 17 119
rect -17 17 17 51
rect -17 -51 17 -17
rect -17 -119 17 -89
rect -17 -187 17 -161
rect -17 -255 17 -233
rect -17 -329 17 -305
rect 201 305 235 329
rect 201 233 235 255
rect 201 161 235 187
rect 201 89 235 119
rect 201 17 235 51
rect 201 -51 235 -17
rect 201 -119 235 -89
rect 201 -187 235 -161
rect 201 -255 235 -233
rect 201 -329 235 -305
rect 315 323 349 357
rect 315 255 349 289
rect 315 187 349 221
rect 315 119 349 153
rect 315 51 349 85
rect 315 -17 349 17
rect 315 -85 349 -51
rect 315 -153 349 -119
rect 315 -221 349 -187
rect 315 -289 349 -255
rect 315 -357 349 -323
rect -349 -465 -315 -391
rect -189 -397 -162 -363
rect -126 -397 -92 -363
rect -56 -397 -29 -363
rect 29 -397 56 -363
rect 92 -397 126 -363
rect 162 -397 189 -363
rect 315 -465 349 -391
rect -349 -499 -221 -465
rect -187 -499 -153 -465
rect -119 -499 -85 -465
rect -51 -499 -17 -465
rect 17 -499 51 -465
rect 85 -499 119 -465
rect 153 -499 187 -465
rect 221 -499 349 -465
<< viali >>
rect -162 363 -160 397
rect -160 363 -128 397
rect -90 363 -58 397
rect -58 363 -56 397
rect 56 363 58 397
rect 58 363 90 397
rect 128 363 160 397
rect 160 363 162 397
rect -235 289 -201 305
rect -235 271 -201 289
rect -235 221 -201 233
rect -235 199 -201 221
rect -235 153 -201 161
rect -235 127 -201 153
rect -235 85 -201 89
rect -235 55 -201 85
rect -235 -17 -201 17
rect -235 -85 -201 -55
rect -235 -89 -201 -85
rect -235 -153 -201 -127
rect -235 -161 -201 -153
rect -235 -221 -201 -199
rect -235 -233 -201 -221
rect -235 -289 -201 -271
rect -235 -305 -201 -289
rect -17 289 17 305
rect -17 271 17 289
rect -17 221 17 233
rect -17 199 17 221
rect -17 153 17 161
rect -17 127 17 153
rect -17 85 17 89
rect -17 55 17 85
rect -17 -17 17 17
rect -17 -85 17 -55
rect -17 -89 17 -85
rect -17 -153 17 -127
rect -17 -161 17 -153
rect -17 -221 17 -199
rect -17 -233 17 -221
rect -17 -289 17 -271
rect -17 -305 17 -289
rect 201 289 235 305
rect 201 271 235 289
rect 201 221 235 233
rect 201 199 235 221
rect 201 153 235 161
rect 201 127 235 153
rect 201 85 235 89
rect 201 55 235 85
rect 201 -17 235 17
rect 201 -85 235 -55
rect 201 -89 235 -85
rect 201 -153 235 -127
rect 201 -161 235 -153
rect 201 -221 235 -199
rect 201 -233 235 -221
rect 201 -289 235 -271
rect 201 -305 235 -289
rect -162 -397 -160 -363
rect -160 -397 -128 -363
rect -90 -397 -58 -363
rect -58 -397 -56 -363
rect 56 -397 58 -363
rect 58 -397 90 -363
rect 128 -397 160 -363
rect 160 -397 162 -363
<< metal1 >>
rect -185 397 -33 403
rect -185 363 -162 397
rect -128 363 -90 397
rect -56 363 -33 397
rect -185 357 -33 363
rect 33 397 185 403
rect 33 363 56 397
rect 90 363 128 397
rect 162 363 185 397
rect 33 357 185 363
rect -241 305 -195 325
rect -241 271 -235 305
rect -201 271 -195 305
rect -241 233 -195 271
rect -241 199 -235 233
rect -201 199 -195 233
rect -241 161 -195 199
rect -241 127 -235 161
rect -201 127 -195 161
rect -241 89 -195 127
rect -241 55 -235 89
rect -201 55 -195 89
rect -241 17 -195 55
rect -241 -17 -235 17
rect -201 -17 -195 17
rect -241 -55 -195 -17
rect -241 -89 -235 -55
rect -201 -89 -195 -55
rect -241 -127 -195 -89
rect -241 -161 -235 -127
rect -201 -161 -195 -127
rect -241 -199 -195 -161
rect -241 -233 -235 -199
rect -201 -233 -195 -199
rect -241 -271 -195 -233
rect -241 -305 -235 -271
rect -201 -305 -195 -271
rect -241 -325 -195 -305
rect -23 305 23 325
rect -23 271 -17 305
rect 17 271 23 305
rect -23 233 23 271
rect -23 199 -17 233
rect 17 199 23 233
rect -23 161 23 199
rect -23 127 -17 161
rect 17 127 23 161
rect -23 89 23 127
rect -23 55 -17 89
rect 17 55 23 89
rect -23 17 23 55
rect -23 -17 -17 17
rect 17 -17 23 17
rect -23 -55 23 -17
rect -23 -89 -17 -55
rect 17 -89 23 -55
rect -23 -127 23 -89
rect -23 -161 -17 -127
rect 17 -161 23 -127
rect -23 -199 23 -161
rect -23 -233 -17 -199
rect 17 -233 23 -199
rect -23 -271 23 -233
rect -23 -305 -17 -271
rect 17 -305 23 -271
rect -23 -325 23 -305
rect 195 305 241 325
rect 195 271 201 305
rect 235 271 241 305
rect 195 233 241 271
rect 195 199 201 233
rect 235 199 241 233
rect 195 161 241 199
rect 195 127 201 161
rect 235 127 241 161
rect 195 89 241 127
rect 195 55 201 89
rect 235 55 241 89
rect 195 17 241 55
rect 195 -17 201 17
rect 235 -17 241 17
rect 195 -55 241 -17
rect 195 -89 201 -55
rect 235 -89 241 -55
rect 195 -127 241 -89
rect 195 -161 201 -127
rect 235 -161 241 -127
rect 195 -199 241 -161
rect 195 -233 201 -199
rect 235 -233 241 -199
rect 195 -271 241 -233
rect 195 -305 201 -271
rect 235 -305 241 -271
rect 195 -325 241 -305
rect -185 -363 -33 -357
rect -185 -397 -162 -363
rect -128 -397 -90 -363
rect -56 -397 -33 -363
rect -185 -403 -33 -397
rect 33 -363 185 -357
rect 33 -397 56 -363
rect 90 -397 128 -363
rect 162 -397 185 -363
rect 33 -403 185 -397
<< properties >>
string FIXED_BBOX -332 -482 332 482
<< end >>
