magic
tech sky130A
magscale 1 2
timestamp 1712737205
<< error_p >>
rect -29 272 29 278
rect -29 238 -17 272
rect -29 232 29 238
rect -29 -238 29 -232
rect -29 -272 -17 -238
rect -29 -278 29 -272
<< pwell >>
rect -216 -400 216 400
<< nmos >>
rect -30 -200 30 200
<< ndiff >>
rect -88 187 -30 200
rect -88 153 -76 187
rect -42 153 -30 187
rect -88 119 -30 153
rect -88 85 -76 119
rect -42 85 -30 119
rect -88 51 -30 85
rect -88 17 -76 51
rect -42 17 -30 51
rect -88 -17 -30 17
rect -88 -51 -76 -17
rect -42 -51 -30 -17
rect -88 -85 -30 -51
rect -88 -119 -76 -85
rect -42 -119 -30 -85
rect -88 -153 -30 -119
rect -88 -187 -76 -153
rect -42 -187 -30 -153
rect -88 -200 -30 -187
rect 30 187 88 200
rect 30 153 42 187
rect 76 153 88 187
rect 30 119 88 153
rect 30 85 42 119
rect 76 85 88 119
rect 30 51 88 85
rect 30 17 42 51
rect 76 17 88 51
rect 30 -17 88 17
rect 30 -51 42 -17
rect 76 -51 88 -17
rect 30 -85 88 -51
rect 30 -119 42 -85
rect 76 -119 88 -85
rect 30 -153 88 -119
rect 30 -187 42 -153
rect 76 -187 88 -153
rect 30 -200 88 -187
<< ndiffc >>
rect -76 153 -42 187
rect -76 85 -42 119
rect -76 17 -42 51
rect -76 -51 -42 -17
rect -76 -119 -42 -85
rect -76 -187 -42 -153
rect 42 153 76 187
rect 42 85 76 119
rect 42 17 76 51
rect 42 -51 76 -17
rect 42 -119 76 -85
rect 42 -187 76 -153
<< psubdiff >>
rect -190 340 -85 374
rect -51 340 -17 374
rect 17 340 51 374
rect 85 340 190 374
rect -190 255 -156 340
rect 156 255 190 340
rect -190 187 -156 221
rect -190 119 -156 153
rect -190 51 -156 85
rect -190 -17 -156 17
rect -190 -85 -156 -51
rect -190 -153 -156 -119
rect -190 -221 -156 -187
rect 156 187 190 221
rect 156 119 190 153
rect 156 51 190 85
rect 156 -17 190 17
rect 156 -85 190 -51
rect 156 -153 190 -119
rect 156 -221 190 -187
rect -190 -340 -156 -255
rect 156 -340 190 -255
rect -190 -374 -85 -340
rect -51 -374 -17 -340
rect 17 -374 51 -340
rect 85 -374 190 -340
<< psubdiffcont >>
rect -85 340 -51 374
rect -17 340 17 374
rect 51 340 85 374
rect -190 221 -156 255
rect 156 221 190 255
rect -190 153 -156 187
rect -190 85 -156 119
rect -190 17 -156 51
rect -190 -51 -156 -17
rect -190 -119 -156 -85
rect -190 -187 -156 -153
rect 156 153 190 187
rect 156 85 190 119
rect 156 17 190 51
rect 156 -51 190 -17
rect 156 -119 190 -85
rect 156 -187 190 -153
rect -190 -255 -156 -221
rect 156 -255 190 -221
rect -85 -374 -51 -340
rect -17 -374 17 -340
rect 51 -374 85 -340
<< poly >>
rect -33 272 33 288
rect -33 238 -17 272
rect 17 238 33 272
rect -33 222 33 238
rect -30 200 30 222
rect -30 -222 30 -200
rect -33 -238 33 -222
rect -33 -272 -17 -238
rect 17 -272 33 -238
rect -33 -288 33 -272
<< polycont >>
rect -17 238 17 272
rect -17 -272 17 -238
<< locali >>
rect -190 340 -85 374
rect -51 340 -17 374
rect 17 340 51 374
rect 85 340 190 374
rect -190 255 -156 340
rect -33 238 -17 272
rect 17 238 33 272
rect 156 255 190 340
rect -190 187 -156 221
rect -190 119 -156 153
rect -190 51 -156 85
rect -190 -17 -156 17
rect -190 -85 -156 -51
rect -190 -153 -156 -119
rect -190 -221 -156 -187
rect -76 187 -42 204
rect -76 119 -42 127
rect -76 51 -42 55
rect -76 -55 -42 -51
rect -76 -127 -42 -119
rect -76 -204 -42 -187
rect 42 187 76 204
rect 42 119 76 127
rect 42 51 76 55
rect 42 -55 76 -51
rect 42 -127 76 -119
rect 42 -204 76 -187
rect 156 187 190 221
rect 156 119 190 153
rect 156 51 190 85
rect 156 -17 190 17
rect 156 -85 190 -51
rect 156 -153 190 -119
rect 156 -221 190 -187
rect -190 -340 -156 -255
rect -33 -272 -17 -238
rect 17 -272 33 -238
rect 156 -340 190 -255
rect -190 -374 -85 -340
rect -51 -374 -17 -340
rect 17 -374 51 -340
rect 85 -374 190 -340
<< viali >>
rect -17 238 17 272
rect -76 153 -42 161
rect -76 127 -42 153
rect -76 85 -42 89
rect -76 55 -42 85
rect -76 -17 -42 17
rect -76 -85 -42 -55
rect -76 -89 -42 -85
rect -76 -153 -42 -127
rect -76 -161 -42 -153
rect 42 153 76 161
rect 42 127 76 153
rect 42 85 76 89
rect 42 55 76 85
rect 42 -17 76 17
rect 42 -85 76 -55
rect 42 -89 76 -85
rect 42 -153 76 -127
rect 42 -161 76 -153
rect -17 -272 17 -238
<< metal1 >>
rect -29 272 29 278
rect -29 238 -17 272
rect 17 238 29 272
rect -29 232 29 238
rect -82 161 -36 200
rect -82 127 -76 161
rect -42 127 -36 161
rect -82 89 -36 127
rect -82 55 -76 89
rect -42 55 -36 89
rect -82 17 -36 55
rect -82 -17 -76 17
rect -42 -17 -36 17
rect -82 -55 -36 -17
rect -82 -89 -76 -55
rect -42 -89 -36 -55
rect -82 -127 -36 -89
rect -82 -161 -76 -127
rect -42 -161 -36 -127
rect -82 -200 -36 -161
rect 36 161 82 200
rect 36 127 42 161
rect 76 127 82 161
rect 36 89 82 127
rect 36 55 42 89
rect 76 55 82 89
rect 36 17 82 55
rect 36 -17 42 17
rect 76 -17 82 17
rect 36 -55 82 -17
rect 36 -89 42 -55
rect 76 -89 82 -55
rect 36 -127 82 -89
rect 36 -161 42 -127
rect 76 -161 82 -127
rect 36 -200 82 -161
rect -29 -238 29 -232
rect -29 -272 -17 -238
rect 17 -272 29 -238
rect -29 -278 29 -272
<< properties >>
string FIXED_BBOX -173 -357 173 357
<< end >>
