magic
tech sky130A
magscale 1 2
timestamp 1712737205
<< nwell >>
rect 3218 152 3338 320
rect 5702 50 5894 318
rect 8164 -2 8440 318
<< pwell >>
rect 3198 -220 3320 -50
rect 5726 -226 5878 -82
rect 8140 -248 8298 -72
<< psubdiff >>
rect 3224 -109 3294 -76
rect 3224 -143 3242 -109
rect 3276 -143 3294 -109
rect 3224 -194 3294 -143
rect 5752 -136 5852 -108
rect 5752 -170 5774 -136
rect 5808 -170 5852 -136
rect 5752 -200 5852 -170
rect 8166 -139 8272 -98
rect 8166 -173 8194 -139
rect 8228 -173 8272 -139
rect 8166 -222 8272 -173
<< nsubdiff >>
rect 3212 254 3298 266
rect 3212 220 3239 254
rect 3273 220 3298 254
rect 3212 192 3298 220
rect 5728 187 5852 262
rect 5728 153 5766 187
rect 5800 153 5852 187
rect 5728 96 5852 153
rect 8222 183 8384 242
rect 8222 149 8288 183
rect 8322 149 8384 183
rect 8222 82 8384 149
<< psubdiffcont >>
rect 3242 -143 3276 -109
rect 5774 -170 5808 -136
rect 8194 -173 8228 -139
<< nsubdiffcont >>
rect 3239 220 3273 254
rect 5766 153 5800 187
rect 8288 149 8322 183
<< locali >>
rect 3116 258 3180 300
rect 3116 254 3292 258
rect 3116 220 3239 254
rect 3273 220 3292 254
rect 3116 206 3292 220
rect 5606 187 5826 204
rect 5606 153 5766 187
rect 5800 153 5826 187
rect 5606 136 5826 153
rect 8064 183 8358 208
rect 8064 149 8288 183
rect 8322 149 8358 183
rect 8064 120 8358 149
rect 3750 50 3816 58
rect 1276 0 1326 18
rect 1276 -34 1284 0
rect 1318 -34 1326 0
rect 3750 16 3766 50
rect 3800 16 3816 50
rect 1276 -52 1326 -34
rect 1526 -34 1568 -24
rect 1526 -68 1530 -34
rect 1564 -68 1568 -34
rect 1526 -78 1568 -68
rect 3036 -30 3070 -8
rect 3750 -22 3816 16
rect 3750 -56 3766 -22
rect 3800 -56 3816 -22
rect 6220 5 6280 38
rect 3750 -64 3816 -56
rect 4006 -39 4062 -28
rect 3036 -86 3070 -64
rect 4006 -73 4017 -39
rect 4051 -73 4062 -39
rect 4006 -84 4062 -73
rect 5522 -38 5556 -26
rect 6220 -29 6233 5
rect 6267 -29 6280 5
rect 6220 -62 6280 -29
rect 6472 -23 6522 -16
rect 6472 -57 6480 -23
rect 6514 -57 6522 -23
rect 6472 -64 6522 -57
rect 7982 -26 8024 -16
rect 7982 -60 7986 -26
rect 8020 -60 8024 -26
rect 7982 -70 8024 -60
rect 5522 -84 5556 -72
rect 3140 -107 3302 -100
rect 3140 -108 3243 -107
rect 3138 -109 3243 -108
rect 2630 -141 2692 -136
rect 2630 -175 2644 -141
rect 2678 -175 2692 -141
rect 3138 -143 3242 -109
rect 3277 -141 3302 -107
rect 3276 -143 3302 -141
rect 3138 -146 3302 -143
rect 3140 -148 3302 -146
rect 5114 -134 5170 -130
rect 5114 -168 5125 -134
rect 5159 -168 5170 -134
rect 5114 -172 5170 -168
rect 5604 -134 5826 -128
rect 5604 -136 5777 -134
rect 5604 -170 5774 -136
rect 5811 -168 5826 -134
rect 5808 -170 5826 -168
rect 2630 -180 2692 -175
rect 5604 -190 5826 -170
rect 7576 -135 7642 -128
rect 7576 -169 7592 -135
rect 7626 -169 7642 -135
rect 7576 -176 7642 -169
rect 8070 -138 8240 -118
rect 8070 -172 8193 -138
rect 8227 -139 8240 -138
rect 8070 -173 8194 -172
rect 8228 -173 8240 -139
rect 8070 -192 8240 -173
<< viali >>
rect 1284 -34 1318 0
rect 3766 16 3800 50
rect 1530 -68 1564 -34
rect 3036 -64 3070 -30
rect 3766 -56 3800 -22
rect 4017 -73 4051 -39
rect 5522 -72 5556 -38
rect 6233 -29 6267 5
rect 6480 -57 6514 -23
rect 7986 -60 8020 -26
rect 3243 -109 3277 -107
rect 2644 -175 2678 -141
rect 3243 -141 3276 -109
rect 3276 -141 3277 -109
rect 5125 -168 5159 -134
rect 5777 -136 5811 -134
rect 5777 -168 5808 -136
rect 5808 -168 5811 -136
rect 7592 -169 7626 -135
rect 8193 -139 8227 -138
rect 8193 -172 8194 -139
rect 8194 -172 8227 -139
<< metal1 >>
rect 2650 440 2850 570
rect 3412 514 3612 630
rect 2650 388 2716 440
rect 2768 388 2850 440
rect 2650 370 2850 388
rect 3410 430 3612 514
rect 5132 449 5332 564
rect 3410 330 3610 430
rect 5132 397 5194 449
rect 5246 397 5332 449
rect 5132 364 5332 397
rect 7608 447 7808 572
rect 7608 395 7643 447
rect 7695 395 7707 447
rect 7759 395 7808 447
rect 7608 372 7808 395
rect 1246 230 5658 330
rect 5664 236 6224 330
rect 974 16 1174 66
rect 3744 50 3822 70
rect 1270 16 1332 30
rect 974 0 1332 16
rect 3744 16 3766 50
rect 3800 16 3822 50
rect 974 -34 1284 0
rect 1318 -34 1332 0
rect 3030 -6 3076 4
rect 3744 -6 3822 16
rect 3030 -10 3822 -6
rect 974 -64 1332 -34
rect 1520 -22 3822 -10
rect 6214 5 6286 50
rect 5516 -16 5562 -14
rect 6214 -16 6233 5
rect 5516 -20 6233 -16
rect 1520 -30 3766 -22
rect 1520 -34 3036 -30
rect 974 -134 1174 -64
rect 1520 -68 1530 -34
rect 1564 -64 3036 -34
rect 3070 -56 3766 -30
rect 3800 -56 3822 -22
rect 3070 -64 3822 -56
rect 1564 -66 3822 -64
rect 1564 -68 3076 -66
rect 1520 -88 3076 -68
rect 3744 -76 3822 -66
rect 3992 -29 6233 -20
rect 6267 -29 6286 5
rect 3992 -38 6286 -29
rect 3992 -39 5522 -38
rect 3992 -73 4017 -39
rect 4051 -72 5522 -39
rect 5556 -66 6286 -38
rect 5556 -72 5562 -66
rect 4051 -73 5562 -72
rect 3992 -86 5562 -73
rect 6214 -74 6286 -66
rect 6460 -16 6534 -10
rect 7976 -16 8030 -4
rect 6460 -23 8030 -16
rect 6460 -57 6480 -23
rect 6514 -26 8030 -23
rect 6514 -57 7986 -26
rect 6460 -60 7986 -57
rect 8020 -60 8030 -26
rect 6460 -70 8030 -60
rect 7976 -82 8030 -70
rect 1520 -90 1574 -88
rect 3030 -98 3076 -88
rect 3994 -90 4074 -86
rect 3214 -107 3306 -94
rect 5516 -96 5562 -86
rect 2618 -132 2790 -130
rect 2618 -141 2716 -132
rect 2618 -175 2644 -141
rect 2678 -175 2716 -141
rect 2618 -184 2716 -175
rect 2768 -184 2790 -132
rect 3214 -141 3243 -107
rect 3277 -141 3306 -107
rect 3214 -154 3306 -141
rect 5102 -125 5276 -124
rect 5102 -134 5198 -125
rect 5102 -168 5125 -134
rect 5159 -168 5198 -134
rect 5102 -177 5198 -168
rect 5250 -177 5276 -125
rect 7564 -126 7752 -122
rect 5760 -134 5828 -126
rect 5760 -168 5777 -134
rect 5811 -168 5828 -134
rect 5760 -176 5828 -168
rect 7564 -135 7671 -126
rect 7564 -169 7592 -135
rect 7626 -169 7671 -135
rect 5102 -178 5276 -177
rect 7564 -178 7671 -169
rect 7723 -178 7752 -126
rect 7564 -182 7752 -178
rect 8178 -138 8242 -110
rect 8178 -172 8193 -138
rect 8227 -172 8242 -138
rect 2618 -186 2790 -184
rect 8178 -200 8242 -172
rect 3180 -310 3756 -212
rect 3392 -528 3618 -310
rect 5654 -318 6214 -224
rect 3406 -588 3606 -528
<< via1 >>
rect 2716 388 2768 440
rect 5194 397 5246 449
rect 7643 395 7695 447
rect 7707 395 7759 447
rect 2716 -184 2768 -132
rect 5198 -177 5250 -125
rect 7671 -178 7723 -126
<< metal2 >>
rect 5186 482 5254 488
rect 2706 460 2778 468
rect 2704 440 2780 460
rect 2704 388 2716 440
rect 2768 388 2780 440
rect 2704 -132 2780 388
rect 2704 -184 2716 -132
rect 2768 -184 2780 -132
rect 2704 -196 2780 -184
rect 5182 449 5254 482
rect 5182 397 5194 449
rect 5246 397 5254 449
rect 5182 -114 5254 397
rect 7638 447 7764 474
rect 7638 395 7643 447
rect 7695 395 7707 447
rect 7759 395 7764 447
rect 7638 368 7764 395
rect 5182 -125 5266 -114
rect 5182 -177 5198 -125
rect 5250 -177 5266 -125
rect 5182 -188 5266 -177
rect 7650 -126 7764 368
rect 7650 -178 7671 -126
rect 7723 -178 7764 -126
rect 7650 -180 7764 -178
rect 7652 -192 7742 -180
use sky130_fd_sc_hd__dfxbp_2  x1
timestamp 1712737205
transform 1 0 1248 0 1 -262
box -38 -48 1970 592
use sky130_fd_sc_hd__dfxbp_2  x2
timestamp 1712737205
transform 1 0 3732 0 1 -262
box -38 -48 1970 592
use sky130_fd_sc_hd__dfxbp_2  x3
timestamp 1712737205
transform 1 0 6196 0 1 -266
box -38 -48 1970 592
<< labels >>
flabel metal1 s 3412 430 3612 630 0 FreeSans 500 0 0 0 VDD
port 1 nsew
flabel metal1 s 3406 -588 3606 -388 0 FreeSans 500 0 0 0 VSS
port 2 nsew
flabel metal1 s 2650 370 2850 570 0 FreeSans 500 0 0 0 Out_2
port 3 nsew
flabel metal1 s 5132 364 5332 564 0 FreeSans 500 0 0 0 Out_4
port 4 nsew
flabel metal1 s 7608 372 7808 572 0 FreeSans 500 0 0 0 Out_8
port 5 nsew
flabel metal1 s 974 -134 1174 66 0 FreeSans 500 0 0 0 Input
port 6 nsew
<< end >>
