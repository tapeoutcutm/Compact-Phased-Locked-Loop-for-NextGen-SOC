magic
tech sky130A
magscale 1 2
timestamp 1712737205
<< error_p >>
rect -88 781 -30 787
rect 30 781 88 787
rect -88 747 -76 781
rect 30 747 42 781
rect -88 741 -30 747
rect 30 741 88 747
rect -88 -747 -30 -741
rect 30 -747 88 -741
rect -88 -781 -76 -747
rect 30 -781 42 -747
rect -88 -787 -30 -781
rect 30 -787 88 -781
<< nwell >>
rect -285 -919 285 919
<< pmos >>
rect -89 -700 -29 700
rect 29 -700 89 700
<< pdiff >>
rect -147 663 -89 700
rect -147 629 -135 663
rect -101 629 -89 663
rect -147 595 -89 629
rect -147 561 -135 595
rect -101 561 -89 595
rect -147 527 -89 561
rect -147 493 -135 527
rect -101 493 -89 527
rect -147 459 -89 493
rect -147 425 -135 459
rect -101 425 -89 459
rect -147 391 -89 425
rect -147 357 -135 391
rect -101 357 -89 391
rect -147 323 -89 357
rect -147 289 -135 323
rect -101 289 -89 323
rect -147 255 -89 289
rect -147 221 -135 255
rect -101 221 -89 255
rect -147 187 -89 221
rect -147 153 -135 187
rect -101 153 -89 187
rect -147 119 -89 153
rect -147 85 -135 119
rect -101 85 -89 119
rect -147 51 -89 85
rect -147 17 -135 51
rect -101 17 -89 51
rect -147 -17 -89 17
rect -147 -51 -135 -17
rect -101 -51 -89 -17
rect -147 -85 -89 -51
rect -147 -119 -135 -85
rect -101 -119 -89 -85
rect -147 -153 -89 -119
rect -147 -187 -135 -153
rect -101 -187 -89 -153
rect -147 -221 -89 -187
rect -147 -255 -135 -221
rect -101 -255 -89 -221
rect -147 -289 -89 -255
rect -147 -323 -135 -289
rect -101 -323 -89 -289
rect -147 -357 -89 -323
rect -147 -391 -135 -357
rect -101 -391 -89 -357
rect -147 -425 -89 -391
rect -147 -459 -135 -425
rect -101 -459 -89 -425
rect -147 -493 -89 -459
rect -147 -527 -135 -493
rect -101 -527 -89 -493
rect -147 -561 -89 -527
rect -147 -595 -135 -561
rect -101 -595 -89 -561
rect -147 -629 -89 -595
rect -147 -663 -135 -629
rect -101 -663 -89 -629
rect -147 -700 -89 -663
rect -29 663 29 700
rect -29 629 -17 663
rect 17 629 29 663
rect -29 595 29 629
rect -29 561 -17 595
rect 17 561 29 595
rect -29 527 29 561
rect -29 493 -17 527
rect 17 493 29 527
rect -29 459 29 493
rect -29 425 -17 459
rect 17 425 29 459
rect -29 391 29 425
rect -29 357 -17 391
rect 17 357 29 391
rect -29 323 29 357
rect -29 289 -17 323
rect 17 289 29 323
rect -29 255 29 289
rect -29 221 -17 255
rect 17 221 29 255
rect -29 187 29 221
rect -29 153 -17 187
rect 17 153 29 187
rect -29 119 29 153
rect -29 85 -17 119
rect 17 85 29 119
rect -29 51 29 85
rect -29 17 -17 51
rect 17 17 29 51
rect -29 -17 29 17
rect -29 -51 -17 -17
rect 17 -51 29 -17
rect -29 -85 29 -51
rect -29 -119 -17 -85
rect 17 -119 29 -85
rect -29 -153 29 -119
rect -29 -187 -17 -153
rect 17 -187 29 -153
rect -29 -221 29 -187
rect -29 -255 -17 -221
rect 17 -255 29 -221
rect -29 -289 29 -255
rect -29 -323 -17 -289
rect 17 -323 29 -289
rect -29 -357 29 -323
rect -29 -391 -17 -357
rect 17 -391 29 -357
rect -29 -425 29 -391
rect -29 -459 -17 -425
rect 17 -459 29 -425
rect -29 -493 29 -459
rect -29 -527 -17 -493
rect 17 -527 29 -493
rect -29 -561 29 -527
rect -29 -595 -17 -561
rect 17 -595 29 -561
rect -29 -629 29 -595
rect -29 -663 -17 -629
rect 17 -663 29 -629
rect -29 -700 29 -663
rect 89 663 147 700
rect 89 629 101 663
rect 135 629 147 663
rect 89 595 147 629
rect 89 561 101 595
rect 135 561 147 595
rect 89 527 147 561
rect 89 493 101 527
rect 135 493 147 527
rect 89 459 147 493
rect 89 425 101 459
rect 135 425 147 459
rect 89 391 147 425
rect 89 357 101 391
rect 135 357 147 391
rect 89 323 147 357
rect 89 289 101 323
rect 135 289 147 323
rect 89 255 147 289
rect 89 221 101 255
rect 135 221 147 255
rect 89 187 147 221
rect 89 153 101 187
rect 135 153 147 187
rect 89 119 147 153
rect 89 85 101 119
rect 135 85 147 119
rect 89 51 147 85
rect 89 17 101 51
rect 135 17 147 51
rect 89 -17 147 17
rect 89 -51 101 -17
rect 135 -51 147 -17
rect 89 -85 147 -51
rect 89 -119 101 -85
rect 135 -119 147 -85
rect 89 -153 147 -119
rect 89 -187 101 -153
rect 135 -187 147 -153
rect 89 -221 147 -187
rect 89 -255 101 -221
rect 135 -255 147 -221
rect 89 -289 147 -255
rect 89 -323 101 -289
rect 135 -323 147 -289
rect 89 -357 147 -323
rect 89 -391 101 -357
rect 135 -391 147 -357
rect 89 -425 147 -391
rect 89 -459 101 -425
rect 135 -459 147 -425
rect 89 -493 147 -459
rect 89 -527 101 -493
rect 135 -527 147 -493
rect 89 -561 147 -527
rect 89 -595 101 -561
rect 135 -595 147 -561
rect 89 -629 147 -595
rect 89 -663 101 -629
rect 135 -663 147 -629
rect 89 -700 147 -663
<< pdiffc >>
rect -135 629 -101 663
rect -135 561 -101 595
rect -135 493 -101 527
rect -135 425 -101 459
rect -135 357 -101 391
rect -135 289 -101 323
rect -135 221 -101 255
rect -135 153 -101 187
rect -135 85 -101 119
rect -135 17 -101 51
rect -135 -51 -101 -17
rect -135 -119 -101 -85
rect -135 -187 -101 -153
rect -135 -255 -101 -221
rect -135 -323 -101 -289
rect -135 -391 -101 -357
rect -135 -459 -101 -425
rect -135 -527 -101 -493
rect -135 -595 -101 -561
rect -135 -663 -101 -629
rect -17 629 17 663
rect -17 561 17 595
rect -17 493 17 527
rect -17 425 17 459
rect -17 357 17 391
rect -17 289 17 323
rect -17 221 17 255
rect -17 153 17 187
rect -17 85 17 119
rect -17 17 17 51
rect -17 -51 17 -17
rect -17 -119 17 -85
rect -17 -187 17 -153
rect -17 -255 17 -221
rect -17 -323 17 -289
rect -17 -391 17 -357
rect -17 -459 17 -425
rect -17 -527 17 -493
rect -17 -595 17 -561
rect -17 -663 17 -629
rect 101 629 135 663
rect 101 561 135 595
rect 101 493 135 527
rect 101 425 135 459
rect 101 357 135 391
rect 101 289 135 323
rect 101 221 135 255
rect 101 153 135 187
rect 101 85 135 119
rect 101 17 135 51
rect 101 -51 135 -17
rect 101 -119 135 -85
rect 101 -187 135 -153
rect 101 -255 135 -221
rect 101 -323 135 -289
rect 101 -391 135 -357
rect 101 -459 135 -425
rect 101 -527 135 -493
rect 101 -595 135 -561
rect 101 -663 135 -629
<< nsubdiff >>
rect -249 849 -153 883
rect -119 849 -85 883
rect -51 849 -17 883
rect 17 849 51 883
rect 85 849 119 883
rect 153 849 249 883
rect -249 765 -215 849
rect 215 765 249 849
rect -249 697 -215 731
rect -249 629 -215 663
rect -249 561 -215 595
rect -249 493 -215 527
rect -249 425 -215 459
rect -249 357 -215 391
rect -249 289 -215 323
rect -249 221 -215 255
rect -249 153 -215 187
rect -249 85 -215 119
rect -249 17 -215 51
rect -249 -51 -215 -17
rect -249 -119 -215 -85
rect -249 -187 -215 -153
rect -249 -255 -215 -221
rect -249 -323 -215 -289
rect -249 -391 -215 -357
rect -249 -459 -215 -425
rect -249 -527 -215 -493
rect -249 -595 -215 -561
rect -249 -663 -215 -629
rect -249 -731 -215 -697
rect 215 697 249 731
rect 215 629 249 663
rect 215 561 249 595
rect 215 493 249 527
rect 215 425 249 459
rect 215 357 249 391
rect 215 289 249 323
rect 215 221 249 255
rect 215 153 249 187
rect 215 85 249 119
rect 215 17 249 51
rect 215 -51 249 -17
rect 215 -119 249 -85
rect 215 -187 249 -153
rect 215 -255 249 -221
rect 215 -323 249 -289
rect 215 -391 249 -357
rect 215 -459 249 -425
rect 215 -527 249 -493
rect 215 -595 249 -561
rect 215 -663 249 -629
rect 215 -731 249 -697
rect -249 -849 -215 -765
rect 215 -849 249 -765
rect -249 -883 -153 -849
rect -119 -883 -85 -849
rect -51 -883 -17 -849
rect 17 -883 51 -849
rect 85 -883 119 -849
rect 153 -883 249 -849
<< nsubdiffcont >>
rect -153 849 -119 883
rect -85 849 -51 883
rect -17 849 17 883
rect 51 849 85 883
rect 119 849 153 883
rect -249 731 -215 765
rect 215 731 249 765
rect -249 663 -215 697
rect -249 595 -215 629
rect -249 527 -215 561
rect -249 459 -215 493
rect -249 391 -215 425
rect -249 323 -215 357
rect -249 255 -215 289
rect -249 187 -215 221
rect -249 119 -215 153
rect -249 51 -215 85
rect -249 -17 -215 17
rect -249 -85 -215 -51
rect -249 -153 -215 -119
rect -249 -221 -215 -187
rect -249 -289 -215 -255
rect -249 -357 -215 -323
rect -249 -425 -215 -391
rect -249 -493 -215 -459
rect -249 -561 -215 -527
rect -249 -629 -215 -595
rect -249 -697 -215 -663
rect 215 663 249 697
rect 215 595 249 629
rect 215 527 249 561
rect 215 459 249 493
rect 215 391 249 425
rect 215 323 249 357
rect 215 255 249 289
rect 215 187 249 221
rect 215 119 249 153
rect 215 51 249 85
rect 215 -17 249 17
rect 215 -85 249 -51
rect 215 -153 249 -119
rect 215 -221 249 -187
rect 215 -289 249 -255
rect 215 -357 249 -323
rect 215 -425 249 -391
rect 215 -493 249 -459
rect 215 -561 249 -527
rect 215 -629 249 -595
rect 215 -697 249 -663
rect -249 -765 -215 -731
rect 215 -765 249 -731
rect -153 -883 -119 -849
rect -85 -883 -51 -849
rect -17 -883 17 -849
rect 51 -883 85 -849
rect 119 -883 153 -849
<< poly >>
rect -92 781 -26 797
rect -92 747 -76 781
rect -42 747 -26 781
rect -92 731 -26 747
rect 26 781 92 797
rect 26 747 42 781
rect 76 747 92 781
rect 26 731 92 747
rect -89 700 -29 731
rect 29 700 89 731
rect -89 -731 -29 -700
rect 29 -731 89 -700
rect -92 -747 -26 -731
rect -92 -781 -76 -747
rect -42 -781 -26 -747
rect -92 -797 -26 -781
rect 26 -747 92 -731
rect 26 -781 42 -747
rect 76 -781 92 -747
rect 26 -797 92 -781
<< polycont >>
rect -76 747 -42 781
rect 42 747 76 781
rect -76 -781 -42 -747
rect 42 -781 76 -747
<< locali >>
rect -249 849 -153 883
rect -119 849 -85 883
rect -51 849 -17 883
rect 17 849 51 883
rect 85 849 119 883
rect 153 849 249 883
rect -249 765 -215 849
rect -92 747 -76 781
rect -42 747 -26 781
rect 26 747 42 781
rect 76 747 92 781
rect 215 765 249 849
rect -249 697 -215 731
rect -249 629 -215 663
rect -249 561 -215 595
rect -249 493 -215 527
rect -249 425 -215 459
rect -249 357 -215 391
rect -249 289 -215 323
rect -249 221 -215 255
rect -249 153 -215 187
rect -249 85 -215 119
rect -249 17 -215 51
rect -249 -51 -215 -17
rect -249 -119 -215 -85
rect -249 -187 -215 -153
rect -249 -255 -215 -221
rect -249 -323 -215 -289
rect -249 -391 -215 -357
rect -249 -459 -215 -425
rect -249 -527 -215 -493
rect -249 -595 -215 -561
rect -249 -663 -215 -629
rect -249 -731 -215 -697
rect -135 665 -101 704
rect -135 595 -101 629
rect -135 527 -101 559
rect -135 459 -101 487
rect -135 391 -101 415
rect -135 323 -101 343
rect -135 255 -101 271
rect -135 187 -101 199
rect -135 119 -101 127
rect -135 51 -101 55
rect -135 -55 -101 -51
rect -135 -127 -101 -119
rect -135 -199 -101 -187
rect -135 -271 -101 -255
rect -135 -343 -101 -323
rect -135 -415 -101 -391
rect -135 -487 -101 -459
rect -135 -559 -101 -527
rect -135 -629 -101 -595
rect -135 -704 -101 -665
rect -17 665 17 704
rect -17 595 17 629
rect -17 527 17 559
rect -17 459 17 487
rect -17 391 17 415
rect -17 323 17 343
rect -17 255 17 271
rect -17 187 17 199
rect -17 119 17 127
rect -17 51 17 55
rect -17 -55 17 -51
rect -17 -127 17 -119
rect -17 -199 17 -187
rect -17 -271 17 -255
rect -17 -343 17 -323
rect -17 -415 17 -391
rect -17 -487 17 -459
rect -17 -559 17 -527
rect -17 -629 17 -595
rect -17 -704 17 -665
rect 101 665 135 704
rect 101 595 135 629
rect 101 527 135 559
rect 101 459 135 487
rect 101 391 135 415
rect 101 323 135 343
rect 101 255 135 271
rect 101 187 135 199
rect 101 119 135 127
rect 101 51 135 55
rect 101 -55 135 -51
rect 101 -127 135 -119
rect 101 -199 135 -187
rect 101 -271 135 -255
rect 101 -343 135 -323
rect 101 -415 135 -391
rect 101 -487 135 -459
rect 101 -559 135 -527
rect 101 -629 135 -595
rect 101 -704 135 -665
rect 215 697 249 731
rect 215 629 249 663
rect 215 561 249 595
rect 215 493 249 527
rect 215 425 249 459
rect 215 357 249 391
rect 215 289 249 323
rect 215 221 249 255
rect 215 153 249 187
rect 215 85 249 119
rect 215 17 249 51
rect 215 -51 249 -17
rect 215 -119 249 -85
rect 215 -187 249 -153
rect 215 -255 249 -221
rect 215 -323 249 -289
rect 215 -391 249 -357
rect 215 -459 249 -425
rect 215 -527 249 -493
rect 215 -595 249 -561
rect 215 -663 249 -629
rect 215 -731 249 -697
rect -249 -849 -215 -765
rect -92 -781 -76 -747
rect -42 -781 -26 -747
rect 26 -781 42 -747
rect 76 -781 92 -747
rect 215 -849 249 -765
rect -249 -883 -153 -849
rect -119 -883 -85 -849
rect -51 -883 -17 -849
rect 17 -883 51 -849
rect 85 -883 119 -849
rect 153 -883 249 -849
<< viali >>
rect -76 747 -42 781
rect 42 747 76 781
rect -135 663 -101 665
rect -135 631 -101 663
rect -135 561 -101 593
rect -135 559 -101 561
rect -135 493 -101 521
rect -135 487 -101 493
rect -135 425 -101 449
rect -135 415 -101 425
rect -135 357 -101 377
rect -135 343 -101 357
rect -135 289 -101 305
rect -135 271 -101 289
rect -135 221 -101 233
rect -135 199 -101 221
rect -135 153 -101 161
rect -135 127 -101 153
rect -135 85 -101 89
rect -135 55 -101 85
rect -135 -17 -101 17
rect -135 -85 -101 -55
rect -135 -89 -101 -85
rect -135 -153 -101 -127
rect -135 -161 -101 -153
rect -135 -221 -101 -199
rect -135 -233 -101 -221
rect -135 -289 -101 -271
rect -135 -305 -101 -289
rect -135 -357 -101 -343
rect -135 -377 -101 -357
rect -135 -425 -101 -415
rect -135 -449 -101 -425
rect -135 -493 -101 -487
rect -135 -521 -101 -493
rect -135 -561 -101 -559
rect -135 -593 -101 -561
rect -135 -663 -101 -631
rect -135 -665 -101 -663
rect -17 663 17 665
rect -17 631 17 663
rect -17 561 17 593
rect -17 559 17 561
rect -17 493 17 521
rect -17 487 17 493
rect -17 425 17 449
rect -17 415 17 425
rect -17 357 17 377
rect -17 343 17 357
rect -17 289 17 305
rect -17 271 17 289
rect -17 221 17 233
rect -17 199 17 221
rect -17 153 17 161
rect -17 127 17 153
rect -17 85 17 89
rect -17 55 17 85
rect -17 -17 17 17
rect -17 -85 17 -55
rect -17 -89 17 -85
rect -17 -153 17 -127
rect -17 -161 17 -153
rect -17 -221 17 -199
rect -17 -233 17 -221
rect -17 -289 17 -271
rect -17 -305 17 -289
rect -17 -357 17 -343
rect -17 -377 17 -357
rect -17 -425 17 -415
rect -17 -449 17 -425
rect -17 -493 17 -487
rect -17 -521 17 -493
rect -17 -561 17 -559
rect -17 -593 17 -561
rect -17 -663 17 -631
rect -17 -665 17 -663
rect 101 663 135 665
rect 101 631 135 663
rect 101 561 135 593
rect 101 559 135 561
rect 101 493 135 521
rect 101 487 135 493
rect 101 425 135 449
rect 101 415 135 425
rect 101 357 135 377
rect 101 343 135 357
rect 101 289 135 305
rect 101 271 135 289
rect 101 221 135 233
rect 101 199 135 221
rect 101 153 135 161
rect 101 127 135 153
rect 101 85 135 89
rect 101 55 135 85
rect 101 -17 135 17
rect 101 -85 135 -55
rect 101 -89 135 -85
rect 101 -153 135 -127
rect 101 -161 135 -153
rect 101 -221 135 -199
rect 101 -233 135 -221
rect 101 -289 135 -271
rect 101 -305 135 -289
rect 101 -357 135 -343
rect 101 -377 135 -357
rect 101 -425 135 -415
rect 101 -449 135 -425
rect 101 -493 135 -487
rect 101 -521 135 -493
rect 101 -561 135 -559
rect 101 -593 135 -561
rect 101 -663 135 -631
rect 101 -665 135 -663
rect -76 -781 -42 -747
rect 42 -781 76 -747
<< metal1 >>
rect -88 781 -30 787
rect -88 747 -76 781
rect -42 747 -30 781
rect -88 741 -30 747
rect 30 781 88 787
rect 30 747 42 781
rect 76 747 88 781
rect 30 741 88 747
rect -141 665 -95 700
rect -141 631 -135 665
rect -101 631 -95 665
rect -141 593 -95 631
rect -141 559 -135 593
rect -101 559 -95 593
rect -141 521 -95 559
rect -141 487 -135 521
rect -101 487 -95 521
rect -141 449 -95 487
rect -141 415 -135 449
rect -101 415 -95 449
rect -141 377 -95 415
rect -141 343 -135 377
rect -101 343 -95 377
rect -141 305 -95 343
rect -141 271 -135 305
rect -101 271 -95 305
rect -141 233 -95 271
rect -141 199 -135 233
rect -101 199 -95 233
rect -141 161 -95 199
rect -141 127 -135 161
rect -101 127 -95 161
rect -141 89 -95 127
rect -141 55 -135 89
rect -101 55 -95 89
rect -141 17 -95 55
rect -141 -17 -135 17
rect -101 -17 -95 17
rect -141 -55 -95 -17
rect -141 -89 -135 -55
rect -101 -89 -95 -55
rect -141 -127 -95 -89
rect -141 -161 -135 -127
rect -101 -161 -95 -127
rect -141 -199 -95 -161
rect -141 -233 -135 -199
rect -101 -233 -95 -199
rect -141 -271 -95 -233
rect -141 -305 -135 -271
rect -101 -305 -95 -271
rect -141 -343 -95 -305
rect -141 -377 -135 -343
rect -101 -377 -95 -343
rect -141 -415 -95 -377
rect -141 -449 -135 -415
rect -101 -449 -95 -415
rect -141 -487 -95 -449
rect -141 -521 -135 -487
rect -101 -521 -95 -487
rect -141 -559 -95 -521
rect -141 -593 -135 -559
rect -101 -593 -95 -559
rect -141 -631 -95 -593
rect -141 -665 -135 -631
rect -101 -665 -95 -631
rect -141 -700 -95 -665
rect -23 665 23 700
rect -23 631 -17 665
rect 17 631 23 665
rect -23 593 23 631
rect -23 559 -17 593
rect 17 559 23 593
rect -23 521 23 559
rect -23 487 -17 521
rect 17 487 23 521
rect -23 449 23 487
rect -23 415 -17 449
rect 17 415 23 449
rect -23 377 23 415
rect -23 343 -17 377
rect 17 343 23 377
rect -23 305 23 343
rect -23 271 -17 305
rect 17 271 23 305
rect -23 233 23 271
rect -23 199 -17 233
rect 17 199 23 233
rect -23 161 23 199
rect -23 127 -17 161
rect 17 127 23 161
rect -23 89 23 127
rect -23 55 -17 89
rect 17 55 23 89
rect -23 17 23 55
rect -23 -17 -17 17
rect 17 -17 23 17
rect -23 -55 23 -17
rect -23 -89 -17 -55
rect 17 -89 23 -55
rect -23 -127 23 -89
rect -23 -161 -17 -127
rect 17 -161 23 -127
rect -23 -199 23 -161
rect -23 -233 -17 -199
rect 17 -233 23 -199
rect -23 -271 23 -233
rect -23 -305 -17 -271
rect 17 -305 23 -271
rect -23 -343 23 -305
rect -23 -377 -17 -343
rect 17 -377 23 -343
rect -23 -415 23 -377
rect -23 -449 -17 -415
rect 17 -449 23 -415
rect -23 -487 23 -449
rect -23 -521 -17 -487
rect 17 -521 23 -487
rect -23 -559 23 -521
rect -23 -593 -17 -559
rect 17 -593 23 -559
rect -23 -631 23 -593
rect -23 -665 -17 -631
rect 17 -665 23 -631
rect -23 -700 23 -665
rect 95 665 141 700
rect 95 631 101 665
rect 135 631 141 665
rect 95 593 141 631
rect 95 559 101 593
rect 135 559 141 593
rect 95 521 141 559
rect 95 487 101 521
rect 135 487 141 521
rect 95 449 141 487
rect 95 415 101 449
rect 135 415 141 449
rect 95 377 141 415
rect 95 343 101 377
rect 135 343 141 377
rect 95 305 141 343
rect 95 271 101 305
rect 135 271 141 305
rect 95 233 141 271
rect 95 199 101 233
rect 135 199 141 233
rect 95 161 141 199
rect 95 127 101 161
rect 135 127 141 161
rect 95 89 141 127
rect 95 55 101 89
rect 135 55 141 89
rect 95 17 141 55
rect 95 -17 101 17
rect 135 -17 141 17
rect 95 -55 141 -17
rect 95 -89 101 -55
rect 135 -89 141 -55
rect 95 -127 141 -89
rect 95 -161 101 -127
rect 135 -161 141 -127
rect 95 -199 141 -161
rect 95 -233 101 -199
rect 135 -233 141 -199
rect 95 -271 141 -233
rect 95 -305 101 -271
rect 135 -305 141 -271
rect 95 -343 141 -305
rect 95 -377 101 -343
rect 135 -377 141 -343
rect 95 -415 141 -377
rect 95 -449 101 -415
rect 135 -449 141 -415
rect 95 -487 141 -449
rect 95 -521 101 -487
rect 135 -521 141 -487
rect 95 -559 141 -521
rect 95 -593 101 -559
rect 135 -593 141 -559
rect 95 -631 141 -593
rect 95 -665 101 -631
rect 135 -665 141 -631
rect 95 -700 141 -665
rect -88 -747 -30 -741
rect -88 -781 -76 -747
rect -42 -781 -30 -747
rect -88 -787 -30 -781
rect 30 -747 88 -741
rect 30 -781 42 -747
rect 76 -781 88 -747
rect 30 -787 88 -781
<< properties >>
string FIXED_BBOX -232 -866 232 866
<< end >>
