VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_vks_pll
  CLASS BLOCK ;
  FOREIGN tt_um_vks_pll ;
  ORIGIN 0.000 0.000 ;
  SIZE 161.000 BY 225.760 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 154.870 224.760 155.170 225.760 ;
    END
  END clk
  PIN ena
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 158.550 224.760 158.850 225.760 ;
    END
  END ena
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 151.190 224.760 151.490 225.760 ;
    END
  END rst_n
  PIN ua[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 5.400000 ;
    PORT
      LAYER li1 ;
        RECT 139.815 26.910 140.145 27.080 ;
        RECT 140.405 26.910 140.735 27.080 ;
        RECT 140.995 26.910 141.325 27.080 ;
        RECT 139.815 20.270 140.145 20.440 ;
        RECT 140.405 20.270 140.735 20.440 ;
        RECT 140.995 20.270 141.325 20.440 ;
      LAYER met1 ;
        RECT 138.420 27.250 141.370 27.280 ;
        RECT 138.070 26.900 141.370 27.250 ;
        RECT 138.070 24.480 138.840 26.900 ;
        RECT 139.835 26.880 140.125 26.900 ;
        RECT 140.425 26.880 140.715 26.900 ;
        RECT 141.015 26.880 141.305 26.900 ;
        RECT 136.790 23.010 138.840 24.480 ;
        RECT 138.070 20.490 138.840 23.010 ;
        RECT 138.070 20.470 141.220 20.490 ;
        RECT 138.070 20.240 141.305 20.470 ;
        RECT 138.130 20.140 141.220 20.240 ;
      LAYER met2 ;
        RECT 136.840 22.960 138.210 24.530 ;
      LAYER met3 ;
        RECT 136.790 22.985 138.260 24.505 ;
      LAYER met4 ;
        RECT 136.835 24.040 138.215 24.485 ;
        RECT 134.670 23.440 138.215 24.040 ;
        RECT 134.670 8.960 135.270 23.440 ;
        RECT 136.835 23.005 138.215 23.440 ;
        RECT 156.560 8.960 157.160 9.000 ;
        RECT 134.670 8.360 157.200 8.960 ;
        RECT 134.670 8.300 135.270 8.360 ;
        RECT 156.560 0.000 157.160 8.360 ;
    END
  END ua[0]
  PIN ua[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.580000 ;
    PORT
      LAYER li1 ;
        RECT 151.035 15.415 151.205 16.455 ;
        RECT 149.330 11.480 149.500 12.520 ;
      LAYER met1 ;
        RECT 155.620 16.440 155.910 16.500 ;
        RECT 151.005 15.960 151.235 16.435 ;
        RECT 155.620 16.400 157.090 16.440 ;
        RECT 150.830 15.560 151.350 15.960 ;
        RECT 154.640 15.680 157.090 16.400 ;
        RECT 151.005 15.435 151.235 15.560 ;
        RECT 154.500 15.160 157.090 15.680 ;
        RECT 155.620 15.110 157.090 15.160 ;
        RECT 155.620 15.040 155.910 15.110 ;
        RECT 149.300 12.270 149.530 12.500 ;
        RECT 149.140 11.830 149.740 12.270 ;
        RECT 149.300 11.500 149.530 11.830 ;
      LAYER met2 ;
        RECT 150.880 15.880 151.300 16.010 ;
        RECT 150.880 15.510 151.560 15.880 ;
        RECT 154.550 15.610 155.620 15.730 ;
        RECT 150.980 14.700 151.560 15.510 ;
        RECT 154.520 15.110 155.620 15.610 ;
        RECT 150.980 14.560 151.630 14.700 ;
        RECT 154.520 14.560 155.450 15.110 ;
        RECT 155.830 15.060 157.040 16.490 ;
        RECT 149.220 13.960 155.460 14.560 ;
        RECT 149.260 13.540 155.460 13.960 ;
        RECT 149.270 12.320 150.060 13.540 ;
        RECT 149.190 11.890 150.060 12.320 ;
        RECT 149.190 11.780 149.690 11.890 ;
      LAYER met3 ;
        RECT 155.780 15.950 157.090 16.465 ;
        RECT 155.250 15.350 159.120 15.950 ;
        RECT 155.780 15.085 157.090 15.350 ;
        RECT 152.785 5.390 153.375 5.415 ;
        RECT 158.520 5.390 159.120 15.350 ;
        RECT 152.780 4.790 159.120 5.390 ;
        RECT 152.785 4.765 153.375 4.790 ;
      LAYER met4 ;
        RECT 134.480 4.790 153.380 5.390 ;
        RECT 134.480 0.000 135.080 4.790 ;
    END
  END ua[1]
  PIN ua[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 20.799999 ;
    PORT
      LAYER li1 ;
        RECT 122.370 21.680 123.170 21.850 ;
        RECT 123.460 21.680 124.260 21.850 ;
        RECT 122.370 17.880 123.170 18.050 ;
        RECT 123.460 17.880 124.260 18.050 ;
        RECT 105.330 11.520 106.130 11.690 ;
        RECT 106.420 11.520 107.220 11.690 ;
        RECT 111.430 11.520 112.230 11.690 ;
        RECT 112.520 11.520 113.320 11.690 ;
        RECT 117.510 11.540 118.310 11.710 ;
        RECT 118.600 11.540 119.400 11.710 ;
        RECT 105.330 7.720 106.130 7.890 ;
        RECT 106.420 7.720 107.220 7.890 ;
        RECT 111.430 7.720 112.230 7.890 ;
        RECT 112.520 7.720 113.320 7.890 ;
        RECT 117.510 7.740 118.310 7.910 ;
        RECT 118.600 7.740 119.400 7.910 ;
      LAYER met1 ;
        RECT 125.120 21.960 125.530 21.970 ;
        RECT 122.340 21.630 125.530 21.960 ;
        RECT 125.120 19.740 125.530 21.630 ;
        RECT 126.820 19.740 128.480 20.240 ;
        RECT 125.120 18.750 128.480 19.740 ;
        RECT 125.120 18.100 125.530 18.750 ;
        RECT 122.390 17.770 125.530 18.100 ;
        RECT 125.120 17.760 125.530 17.770 ;
        RECT 125.900 18.510 128.480 18.750 ;
        RECT 120.640 11.920 121.140 11.930 ;
        RECT 105.270 11.490 121.140 11.920 ;
        RECT 120.640 10.700 121.140 11.490 ;
        RECT 125.900 10.700 126.860 18.510 ;
        RECT 120.640 9.750 126.860 10.700 ;
        RECT 117.530 7.930 118.290 7.940 ;
        RECT 118.620 7.930 119.380 7.940 ;
        RECT 120.640 7.930 121.140 9.750 ;
        RECT 105.290 7.540 121.140 7.930 ;
        RECT 105.290 7.500 121.110 7.540 ;
      LAYER met2 ;
        RECT 126.870 18.460 128.430 20.290 ;
      LAYER met3 ;
        RECT 126.820 18.485 128.480 20.265 ;
      LAYER met4 ;
        RECT 126.865 18.505 128.435 20.245 ;
        RECT 127.260 4.440 127.860 18.505 ;
        RECT 112.400 3.840 127.860 4.440 ;
        RECT 112.400 0.000 113.000 3.840 ;
    END
  END ua[2]
  PIN ua[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.022500 ;
    PORT
      LAYER li1 ;
        RECT 99.970 18.845 100.140 20.885 ;
        RECT 100.930 18.845 101.100 20.885 ;
        RECT 100.820 13.850 100.990 16.140 ;
      LAYER met1 ;
        RECT 99.940 19.370 100.170 20.865 ;
        RECT 99.870 18.950 100.230 19.370 ;
        RECT 100.900 19.340 101.130 20.865 ;
        RECT 99.940 18.865 100.170 18.950 ;
        RECT 100.840 18.920 101.200 19.340 ;
        RECT 100.900 18.865 101.130 18.920 ;
        RECT 96.580 17.810 98.930 18.150 ;
        RECT 100.670 17.810 101.170 17.830 ;
        RECT 96.580 17.350 101.170 17.810 ;
        RECT 96.580 17.310 101.080 17.350 ;
        RECT 96.580 17.060 98.930 17.310 ;
        RECT 97.770 17.020 98.770 17.060 ;
        RECT 100.790 16.100 101.020 16.120 ;
        RECT 100.740 15.540 101.100 16.100 ;
        RECT 100.790 13.870 101.020 15.540 ;
      LAYER met2 ;
        RECT 99.920 19.360 100.180 19.420 ;
        RECT 100.890 19.360 101.150 19.390 ;
        RECT 99.880 18.930 101.160 19.360 ;
        RECT 99.920 18.900 100.180 18.930 ;
        RECT 100.730 18.870 101.150 18.930 ;
        RECT 96.630 17.010 98.880 18.200 ;
        RECT 100.730 17.880 101.090 18.870 ;
        RECT 100.720 17.300 101.120 17.880 ;
        RECT 100.730 15.540 101.090 17.300 ;
        RECT 100.790 15.490 101.050 15.540 ;
      LAYER met3 ;
        RECT 96.580 17.035 98.930 18.175 ;
      LAYER met4 ;
        RECT 96.625 17.650 98.885 18.155 ;
        RECT 90.320 17.055 98.885 17.650 ;
        RECT 90.320 17.050 98.770 17.055 ;
        RECT 90.320 0.000 90.920 17.050 ;
    END
  END ua[3]
  PIN ua[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 68.240 0.000 68.840 1.000 ;
    END
  END ua[4]
  PIN ua[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 46.160 0.000 46.760 1.000 ;
    END
  END ua[5]
  PIN ua[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 24.080 0.000 24.680 1.000 ;
    END
  END ua[6]
  PIN ua[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 2.000 0.000 2.600 1.000 ;
    END
  END ua[7]
  PIN ui_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.000000 ;
    PORT
      LAYER li1 ;
        RECT 151.265 16.670 153.265 16.840 ;
        RECT 151.265 15.030 153.265 15.200 ;
      LAYER met1 ;
        RECT 148.560 17.130 149.560 17.150 ;
        RECT 148.560 16.870 151.850 17.130 ;
        RECT 148.560 16.700 153.245 16.870 ;
        RECT 147.210 16.470 148.350 16.580 ;
        RECT 148.560 16.470 149.610 16.700 ;
        RECT 151.285 16.640 153.245 16.700 ;
        RECT 147.210 15.760 149.610 16.470 ;
        RECT 147.210 15.420 149.750 15.760 ;
        RECT 148.280 15.360 149.750 15.420 ;
        RECT 148.400 15.350 149.750 15.360 ;
        RECT 148.630 15.280 149.750 15.350 ;
        RECT 148.630 15.230 151.890 15.280 ;
        RECT 148.630 15.000 153.245 15.230 ;
        RECT 148.710 14.880 152.040 15.000 ;
        RECT 148.750 14.860 152.040 14.880 ;
        RECT 151.890 14.670 152.040 14.860 ;
      LAYER met2 ;
        RECT 147.260 15.370 148.300 16.630 ;
      LAYER met3 ;
        RECT 147.210 15.395 148.350 16.605 ;
      LAYER met4 ;
        RECT 147.510 43.330 147.815 225.750 ;
        RECT 147.505 40.195 147.820 43.330 ;
        RECT 147.510 40.185 147.815 40.195 ;
        RECT 147.515 16.585 147.815 40.185 ;
        RECT 147.255 15.415 148.305 16.585 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 5.000000 ;
    PORT
      LAYER li1 ;
        RECT 149.560 12.690 154.560 12.860 ;
        RECT 149.560 11.140 154.560 11.310 ;
      LAYER met1 ;
        RECT 147.360 12.890 150.370 13.120 ;
        RECT 147.360 12.780 154.540 12.890 ;
        RECT 147.270 12.680 154.540 12.780 ;
        RECT 147.270 12.530 148.420 12.680 ;
        RECT 149.580 12.660 154.540 12.680 ;
        RECT 147.270 12.510 148.290 12.530 ;
        RECT 147.290 12.280 148.290 12.510 ;
        RECT 146.930 11.670 148.290 12.280 ;
        RECT 146.930 11.340 148.350 11.670 ;
        RECT 146.930 11.110 154.540 11.340 ;
        RECT 146.930 10.920 150.400 11.110 ;
        RECT 147.390 10.900 150.400 10.920 ;
      LAYER met2 ;
        RECT 146.980 10.870 148.040 12.330 ;
      LAYER met3 ;
        RECT 146.930 10.895 148.090 12.305 ;
      LAYER met4 ;
        RECT 143.830 12.090 144.130 225.760 ;
        RECT 146.975 12.090 148.045 12.285 ;
        RECT 143.830 11.790 148.045 12.090 ;
        RECT 146.975 10.915 148.045 11.790 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER li1 ;
        RECT 134.495 183.160 135.145 183.510 ;
        RECT 134.610 181.790 135.110 183.160 ;
      LAYER met1 ;
        RECT 139.980 219.220 140.680 222.010 ;
        RECT 134.580 182.450 135.140 182.510 ;
        RECT 134.380 182.040 135.380 182.450 ;
        RECT 140.140 182.040 140.480 219.220 ;
        RECT 134.380 181.700 140.480 182.040 ;
        RECT 134.380 181.450 135.380 181.700 ;
      LAYER met2 ;
        RECT 140.030 219.170 140.630 222.060 ;
      LAYER met3 ;
        RECT 139.980 219.195 140.680 222.035 ;
      LAYER met4 ;
        RECT 140.150 222.015 140.450 225.760 ;
        RECT 140.025 219.215 140.635 222.015 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER li1 ;
        RECT 10.510 212.315 10.860 212.965 ;
      LAYER met1 ;
        RECT 7.700 222.130 8.860 222.150 ;
        RECT 6.740 221.310 9.860 222.130 ;
        RECT 7.700 213.140 8.860 221.310 ;
        RECT 7.620 212.910 8.890 213.140 ;
        RECT 7.620 212.580 10.850 212.910 ;
        RECT 7.620 211.980 8.890 212.580 ;
      LAYER met2 ;
        RECT 6.790 221.260 9.810 222.180 ;
      LAYER met3 ;
        RECT 6.740 222.060 9.860 222.155 ;
        RECT 6.660 221.850 9.860 222.060 ;
        RECT 136.110 221.850 136.890 222.130 ;
        RECT 6.660 221.760 136.890 221.850 ;
        RECT 6.740 221.550 136.890 221.760 ;
        RECT 6.740 221.285 9.860 221.550 ;
        RECT 136.110 221.530 136.890 221.550 ;
      LAYER met4 ;
        RECT 136.470 222.075 136.770 225.760 ;
        RECT 136.455 221.745 136.785 222.075 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER li1 ;
        RECT 11.230 200.635 11.580 201.285 ;
      LAYER met1 ;
        RECT 8.000 201.300 8.910 202.790 ;
        RECT 8.000 201.050 10.770 201.300 ;
        RECT 11.250 201.050 11.560 201.120 ;
        RECT 8.000 200.650 11.560 201.050 ;
        RECT 8.000 200.300 10.770 200.650 ;
        RECT 8.000 199.800 9.040 200.300 ;
        RECT 8.040 199.780 9.040 199.800 ;
      LAYER met2 ;
        RECT 81.410 209.910 85.680 210.050 ;
        RECT 8.110 209.610 85.680 209.910 ;
        RECT 8.110 202.840 8.410 209.610 ;
        RECT 81.410 209.520 85.680 209.610 ;
        RECT 8.050 199.750 8.860 202.840 ;
      LAYER met3 ;
        RECT 81.360 209.910 85.730 210.025 ;
        RECT 130.950 209.910 131.760 211.380 ;
        RECT 81.360 209.610 131.770 209.910 ;
        RECT 81.360 209.545 85.730 209.610 ;
      LAYER met4 ;
        RECT 132.790 224.410 133.090 225.760 ;
        RECT 131.160 224.110 133.090 224.410 ;
        RECT 131.160 211.385 131.460 224.110 ;
        RECT 130.995 209.645 131.715 211.385 ;
        RECT 131.160 209.620 131.460 209.645 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 129.110 224.760 129.410 225.760 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 125.430 224.760 125.730 225.760 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 121.750 224.760 122.050 225.760 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER li1 ;
        RECT 115.890 204.730 116.240 204.815 ;
        RECT 115.890 204.170 116.530 204.730 ;
        RECT 115.890 204.165 116.240 204.170 ;
      LAYER met1 ;
        RECT 117.000 204.860 118.430 204.990 ;
        RECT 116.330 204.790 118.430 204.860 ;
        RECT 116.320 204.730 118.430 204.790 ;
        RECT 116.110 204.260 118.430 204.730 ;
        RECT 116.320 204.190 118.430 204.260 ;
        RECT 116.330 203.920 118.430 204.190 ;
        RECT 116.330 203.860 117.330 203.920 ;
      LAYER met2 ;
        RECT 117.050 203.870 118.380 205.040 ;
      LAYER met3 ;
        RECT 117.000 203.895 118.430 205.015 ;
      LAYER met4 ;
        RECT 118.070 204.995 118.370 225.760 ;
        RECT 117.045 203.915 118.385 204.995 ;
        RECT 118.070 203.880 118.370 203.915 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 114.390 224.760 114.690 225.760 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER li1 ;
        RECT 76.400 219.410 76.750 219.415 ;
        RECT 77.030 219.410 77.490 219.510 ;
        RECT 76.400 218.780 77.490 219.410 ;
        RECT 76.400 218.765 76.750 218.780 ;
        RECT 77.030 218.510 77.490 218.780 ;
      LAYER met1 ;
        RECT 77.000 219.410 77.520 219.570 ;
        RECT 76.460 218.770 77.520 219.410 ;
        RECT 77.000 218.450 77.520 218.770 ;
        RECT 79.070 219.460 80.070 219.570 ;
        RECT 79.070 218.920 111.250 219.460 ;
        RECT 79.070 218.570 80.070 218.920 ;
      LAYER met2 ;
        RECT 76.930 219.460 79.210 219.480 ;
        RECT 76.510 219.450 79.210 219.460 ;
        RECT 76.510 218.720 79.610 219.450 ;
        RECT 109.820 218.870 111.200 219.510 ;
        RECT 76.930 218.710 79.610 218.720 ;
      LAYER met3 ;
        RECT 109.770 218.895 111.250 219.485 ;
      LAYER met4 ;
        RECT 110.710 219.465 111.010 225.760 ;
        RECT 109.815 218.915 111.205 219.465 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER li1 ;
        RECT 76.400 212.730 76.750 212.735 ;
        RECT 77.100 212.730 77.620 213.050 ;
        RECT 76.400 212.090 77.620 212.730 ;
        RECT 76.400 212.085 76.750 212.090 ;
        RECT 77.100 211.930 77.620 212.090 ;
      LAYER met1 ;
        RECT 76.980 213.110 77.880 213.200 ;
        RECT 106.380 213.110 108.070 213.810 ;
        RECT 76.980 212.800 108.070 213.110 ;
        RECT 76.430 212.450 108.070 212.800 ;
        RECT 76.430 212.360 77.880 212.450 ;
        RECT 76.430 212.060 77.650 212.360 ;
        RECT 79.020 212.060 80.070 212.450 ;
        RECT 106.380 212.240 108.070 212.450 ;
        RECT 77.070 211.870 77.650 212.060 ;
        RECT 79.070 211.950 80.070 212.060 ;
      LAYER met2 ;
        RECT 77.010 212.850 77.850 213.230 ;
        RECT 76.480 212.010 79.490 212.850 ;
        RECT 106.500 212.270 107.790 213.660 ;
      LAYER met3 ;
        RECT 106.530 212.345 107.720 213.525 ;
      LAYER met4 ;
        RECT 107.030 213.505 107.330 225.760 ;
        RECT 106.575 212.365 107.675 213.505 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 103.350 224.760 103.650 225.760 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 99.670 224.760 99.970 225.760 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER li1 ;
        RECT 107.630 195.350 107.980 195.365 ;
        RECT 107.630 194.750 110.570 195.350 ;
        RECT 107.630 194.715 107.980 194.750 ;
      LAYER met1 ;
        RECT 109.990 195.380 111.680 195.540 ;
        RECT 109.770 194.720 111.680 195.380 ;
        RECT 109.990 194.540 111.680 194.720 ;
        RECT 110.710 194.420 111.680 194.540 ;
      LAYER met2 ;
        RECT 110.760 194.370 111.630 195.590 ;
      LAYER met3 ;
        RECT 95.830 211.810 96.580 211.920 ;
        RECT 119.550 211.810 120.380 211.990 ;
        RECT 95.830 211.510 120.380 211.810 ;
        RECT 95.830 211.270 96.580 211.510 ;
        RECT 119.550 211.270 120.380 211.510 ;
        RECT 110.710 194.395 111.680 195.565 ;
      LAYER met4 ;
        RECT 95.990 211.875 96.290 225.760 ;
        RECT 119.770 211.925 120.070 211.940 ;
        RECT 95.895 211.285 96.455 211.875 ;
        RECT 119.675 211.335 120.235 211.925 ;
        RECT 119.680 211.320 120.210 211.335 ;
        RECT 110.755 195.050 111.635 195.545 ;
        RECT 119.910 195.050 120.210 211.320 ;
        RECT 110.755 194.750 120.240 195.050 ;
        RECT 110.755 194.415 111.635 194.750 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER li1 ;
        RECT 107.510 186.610 107.860 186.615 ;
        RECT 107.510 185.980 110.450 186.610 ;
        RECT 107.510 185.970 109.740 185.980 ;
        RECT 107.510 185.965 107.860 185.970 ;
      LAYER met1 ;
        RECT 110.640 186.800 111.660 186.810 ;
        RECT 109.880 186.640 111.660 186.800 ;
        RECT 109.590 185.950 111.660 186.640 ;
        RECT 109.880 185.800 111.660 185.950 ;
      LAYER met2 ;
        RECT 110.690 185.750 111.610 186.860 ;
      LAYER met3 ;
        RECT 121.000 211.540 121.880 212.210 ;
        RECT 92.140 210.960 93.090 211.300 ;
        RECT 120.960 211.240 121.880 211.540 ;
        RECT 92.140 210.810 93.240 210.960 ;
        RECT 121.000 210.810 121.880 211.240 ;
        RECT 92.140 210.510 121.880 210.810 ;
        RECT 92.140 210.280 93.090 210.510 ;
        RECT 121.000 210.490 121.880 210.510 ;
        RECT 110.640 185.775 111.660 186.835 ;
      LAYER met4 ;
        RECT 92.310 211.265 92.610 225.760 ;
        RECT 92.295 210.345 93.025 211.265 ;
        RECT 121.035 210.515 121.815 212.145 ;
        RECT 110.685 186.460 111.615 186.815 ;
        RECT 121.500 186.460 121.800 210.515 ;
        RECT 110.685 186.160 121.800 186.460 ;
        RECT 110.685 185.795 111.615 186.160 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 67.596802 ;
    PORT
      LAYER pwell ;
        RECT 56.940 217.870 57.620 218.860 ;
        RECT 135.075 215.710 135.985 219.395 ;
        RECT 63.060 214.535 63.740 215.430 ;
        RECT 64.735 215.375 66.325 215.465 ;
        RECT 63.755 214.555 66.325 215.375 ;
        RECT 63.755 214.535 63.895 214.555 ;
        RECT 63.060 214.440 63.895 214.535 ;
        RECT 63.725 214.365 63.895 214.440 ;
        RECT 135.305 214.170 135.985 215.710 ;
        RECT 19.170 212.880 20.080 213.770 ;
        RECT 31.980 212.820 32.890 213.710 ;
        RECT 43.880 212.850 44.790 213.740 ;
        RECT 135.085 213.260 135.985 214.170 ;
        RECT 59.770 211.190 60.450 212.180 ;
        RECT 135.305 210.055 135.985 213.260 ;
        RECT 135.305 209.885 136.175 210.055 ;
        RECT 135.305 209.745 135.985 209.885 ;
        RECT 135.310 205.975 135.880 209.745 ;
        RECT 85.520 203.210 86.270 204.260 ;
        RECT 135.055 202.290 135.965 205.975 ;
        RECT 20.790 200.675 21.530 200.770 ;
        RECT 135.285 200.750 135.965 202.290 ;
        RECT 33.210 200.675 34.520 200.680 ;
        RECT 14.660 200.445 15.570 200.665 ;
        RECT 17.110 200.445 21.530 200.675 ;
        RECT 27.080 200.445 27.990 200.665 ;
        RECT 29.530 200.445 34.520 200.675 ;
        RECT 45.530 200.655 46.380 200.660 ;
        RECT 11.145 199.790 21.530 200.445 ;
        RECT 11.145 199.765 20.795 199.790 ;
        RECT 23.565 199.770 34.520 200.445 ;
        RECT 39.400 200.425 40.310 200.645 ;
        RECT 41.850 200.425 46.380 200.655 ;
        RECT 23.565 199.765 33.215 199.770 ;
        RECT 11.285 199.575 11.455 199.765 ;
        RECT 23.705 199.575 23.875 199.765 ;
        RECT 35.885 199.750 46.380 200.425 ;
        RECT 135.065 199.840 135.965 200.750 ;
        RECT 35.885 199.745 45.535 199.750 ;
        RECT 36.025 199.555 36.195 199.745 ;
        RECT 135.285 196.635 135.965 199.840 ;
        RECT 135.285 196.465 136.155 196.635 ;
        RECT 135.285 196.325 135.965 196.465 ;
        RECT 96.010 194.755 97.660 194.770 ;
        RECT 96.010 194.525 99.420 194.755 ;
        RECT 102.625 194.525 103.555 194.745 ;
        RECT 96.010 193.845 108.065 194.525 ;
        RECT 96.010 193.770 97.660 193.845 ;
        RECT 107.755 193.655 107.925 193.845 ;
        RECT 135.380 192.725 135.950 196.325 ;
        RECT 97.910 190.315 99.070 190.350 ;
        RECT 99.925 190.315 101.515 190.405 ;
        RECT 97.910 189.600 101.515 190.315 ;
        RECT 98.945 189.495 101.515 189.600 ;
        RECT 98.945 189.475 99.085 189.495 ;
        RECT 98.915 189.305 99.085 189.475 ;
        RECT 135.105 189.040 136.015 192.725 ;
        RECT 135.335 187.500 136.015 189.040 ;
        RECT 135.115 186.590 136.015 187.500 ;
        RECT 97.020 185.830 99.300 186.005 ;
        RECT 95.910 185.775 99.300 185.830 ;
        RECT 102.505 185.775 103.435 185.995 ;
        RECT 95.910 185.180 107.945 185.775 ;
        RECT 97.020 185.095 107.945 185.180 ;
        RECT 107.635 184.905 107.805 185.095 ;
        RECT 135.335 183.385 136.015 186.590 ;
        RECT 135.335 183.260 136.205 183.385 ;
        RECT 135.330 183.215 136.205 183.260 ;
        RECT 135.330 182.240 136.060 183.215 ;
        RECT 121.440 17.240 125.190 22.490 ;
        RECT 99.640 12.870 102.170 17.120 ;
        RECT 104.440 12.940 108.090 17.190 ;
        RECT 110.530 12.920 114.180 17.170 ;
        RECT 116.540 12.930 120.190 17.180 ;
        RECT 137.115 14.065 139.275 18.065 ;
        RECT 140.865 14.525 143.025 18.525 ;
        RECT 144.150 13.860 146.510 16.560 ;
        RECT 104.400 7.080 108.150 12.330 ;
        RECT 110.500 7.080 114.250 12.330 ;
        RECT 116.580 7.100 120.330 12.350 ;
        RECT 148.630 10.500 155.490 13.500 ;
      LAYER li1 ;
        RECT 136.005 219.305 136.175 219.400 ;
        RECT 135.185 219.055 136.175 219.305 ;
        RECT 57.070 217.900 57.490 218.730 ;
        RECT 57.905 217.900 58.155 218.340 ;
        RECT 57.070 217.875 58.155 217.900 ;
        RECT 58.825 217.875 58.995 218.335 ;
        RECT 59.665 217.875 59.930 218.335 ;
        RECT 60.585 217.875 60.835 218.340 ;
        RECT 61.505 217.875 61.675 218.335 ;
        RECT 62.345 217.875 62.610 218.335 ;
        RECT 63.265 217.875 63.515 218.340 ;
        RECT 64.185 217.875 64.355 218.335 ;
        RECT 65.025 217.875 65.290 218.335 ;
        RECT 66.080 217.875 66.250 218.720 ;
        RECT 66.970 217.875 67.140 218.615 ;
        RECT 136.005 218.460 136.175 219.055 ;
        RECT 67.850 217.875 68.085 218.335 ;
        RECT 69.945 217.875 70.135 218.315 ;
        RECT 72.035 217.875 72.365 218.335 ;
        RECT 74.965 217.875 75.295 218.235 ;
        RECT 75.995 217.875 76.325 218.255 ;
        RECT 135.265 218.130 136.175 218.460 ;
        RECT 57.070 217.710 60.060 217.875 ;
        RECT 57.760 217.705 60.060 217.710 ;
        RECT 60.440 217.705 62.740 217.875 ;
        RECT 63.120 217.705 65.420 217.875 ;
        RECT 65.800 217.705 76.840 217.875 ;
        RECT 136.005 217.310 136.175 218.130 ;
        RECT 135.490 217.140 136.175 217.310 ;
        RECT 136.005 216.470 136.175 217.140 ;
        RECT 135.395 216.300 136.175 216.470 ;
        RECT 136.005 215.535 136.175 216.300 ;
        RECT 63.190 214.540 63.610 215.300 ;
        RECT 64.825 214.540 65.075 214.995 ;
        RECT 63.190 214.535 65.075 214.540 ;
        RECT 65.965 214.535 66.255 215.335 ;
        RECT 135.475 215.325 136.175 215.535 ;
        RECT 66.850 214.535 67.115 214.995 ;
        RECT 67.785 214.535 67.955 214.995 ;
        RECT 68.625 214.535 68.875 215.000 ;
        RECT 63.190 214.370 66.340 214.535 ;
        RECT 63.580 214.365 66.340 214.370 ;
        RECT 66.720 214.365 69.020 214.535 ;
        RECT 10.420 213.855 19.160 214.025 ;
        RECT 23.220 213.865 31.960 214.035 ;
        RECT 35.130 213.865 43.870 214.035 ;
        RECT 10.935 213.475 11.265 213.855 ;
        RECT 11.875 213.395 12.125 213.855 ;
        RECT 13.820 213.355 14.190 213.855 ;
        RECT 16.005 213.325 16.215 213.855 ;
        RECT 16.980 213.245 17.150 213.855 ;
        RECT 18.325 213.395 18.645 213.855 ;
        RECT 19.330 213.040 19.910 213.620 ;
        RECT 23.735 213.485 24.065 213.865 ;
        RECT 24.675 213.405 24.925 213.865 ;
        RECT 26.620 213.365 26.990 213.865 ;
        RECT 28.805 213.335 29.015 213.865 ;
        RECT 29.780 213.255 29.950 213.865 ;
        RECT 31.125 213.405 31.445 213.865 ;
        RECT 32.140 212.980 32.720 213.560 ;
        RECT 35.645 213.485 35.975 213.865 ;
        RECT 36.585 213.405 36.835 213.865 ;
        RECT 38.530 213.365 38.900 213.865 ;
        RECT 40.715 213.335 40.925 213.865 ;
        RECT 41.690 213.255 41.860 213.865 ;
        RECT 43.035 213.405 43.355 213.865 ;
        RECT 44.040 213.010 44.620 213.590 ;
        RECT 136.005 213.510 136.175 215.325 ;
        RECT 135.505 213.140 136.175 213.510 ;
        RECT 59.900 211.210 60.320 212.050 ;
        RECT 60.775 211.210 61.025 211.660 ;
        RECT 59.900 211.195 61.025 211.210 ;
        RECT 61.695 211.195 61.865 211.655 ;
        RECT 62.535 211.195 62.800 211.655 ;
        RECT 63.455 211.195 63.705 211.660 ;
        RECT 64.375 211.195 64.545 211.655 ;
        RECT 65.215 211.195 65.480 211.655 ;
        RECT 66.080 211.195 66.250 212.040 ;
        RECT 66.970 211.195 67.140 211.935 ;
        RECT 67.850 211.195 68.085 211.655 ;
        RECT 69.945 211.195 70.135 211.635 ;
        RECT 72.035 211.195 72.365 211.655 ;
        RECT 74.965 211.195 75.295 211.555 ;
        RECT 75.995 211.195 76.325 211.575 ;
        RECT 136.005 211.445 136.175 213.140 ;
        RECT 135.545 211.195 136.175 211.445 ;
        RECT 59.900 211.030 62.930 211.195 ;
        RECT 60.630 211.025 62.930 211.030 ;
        RECT 63.310 211.025 65.610 211.195 ;
        RECT 65.800 211.025 76.840 211.195 ;
        RECT 136.005 210.585 136.175 211.195 ;
        RECT 135.625 210.255 136.175 210.585 ;
        RECT 136.005 209.740 136.175 210.255 ;
        RECT 135.985 205.885 136.155 205.980 ;
        RECT 135.165 205.635 136.155 205.885 ;
        RECT 135.985 205.040 136.155 205.635 ;
        RECT 135.245 204.710 136.155 205.040 ;
        RECT 85.650 203.340 86.140 204.130 ;
        RECT 86.735 203.340 86.945 204.095 ;
        RECT 85.650 203.275 86.945 203.340 ;
        RECT 87.615 203.275 87.845 204.095 ;
        RECT 88.305 203.275 88.515 204.095 ;
        RECT 89.185 203.275 89.415 204.095 ;
        RECT 135.985 203.890 136.155 204.710 ;
        RECT 90.285 203.275 90.605 203.735 ;
        RECT 91.780 203.275 91.950 203.885 ;
        RECT 92.715 203.275 92.925 203.805 ;
        RECT 94.740 203.275 95.110 203.775 ;
        RECT 96.805 203.275 97.055 203.735 ;
        RECT 97.665 203.275 97.995 203.655 ;
        RECT 99.195 203.275 99.515 203.735 ;
        RECT 100.690 203.275 100.860 203.885 ;
        RECT 101.625 203.275 101.835 203.805 ;
        RECT 103.650 203.275 104.020 203.775 ;
        RECT 105.715 203.275 105.965 203.735 ;
        RECT 106.575 203.275 106.905 203.655 ;
        RECT 108.105 203.275 108.425 203.735 ;
        RECT 109.600 203.275 109.770 203.885 ;
        RECT 110.535 203.275 110.745 203.805 ;
        RECT 112.560 203.275 112.930 203.775 ;
        RECT 114.625 203.275 114.875 203.735 ;
        RECT 135.470 203.720 136.155 203.890 ;
        RECT 115.485 203.275 115.815 203.655 ;
        RECT 85.650 203.110 87.970 203.275 ;
        RECT 86.590 203.105 87.970 203.110 ;
        RECT 88.160 203.105 89.540 203.275 ;
        RECT 89.770 203.105 98.510 203.275 ;
        RECT 98.680 203.105 107.420 203.275 ;
        RECT 107.590 203.105 116.330 203.275 ;
        RECT 135.985 203.050 136.155 203.720 ;
        RECT 135.375 202.880 136.155 203.050 ;
        RECT 135.985 202.115 136.155 202.880 ;
        RECT 135.455 201.905 136.155 202.115 ;
        RECT 11.655 199.745 11.985 200.125 ;
        RECT 12.595 199.745 12.845 200.205 ;
        RECT 14.540 199.745 14.910 200.245 ;
        RECT 16.725 199.745 16.935 200.275 ;
        RECT 17.700 199.745 17.870 200.355 ;
        RECT 18.540 199.745 18.710 200.260 ;
        RECT 19.530 199.745 19.860 200.485 ;
        RECT 20.455 200.470 20.705 200.565 ;
        RECT 20.455 200.230 21.410 200.470 ;
        RECT 20.455 199.745 20.705 200.230 ;
        RECT 24.075 199.745 24.405 200.125 ;
        RECT 25.015 199.745 25.265 200.205 ;
        RECT 26.960 199.745 27.330 200.245 ;
        RECT 29.145 199.745 29.355 200.275 ;
        RECT 30.120 199.745 30.290 200.355 ;
        RECT 30.960 199.745 31.130 200.260 ;
        RECT 31.950 199.745 32.280 200.485 ;
        RECT 32.875 200.330 33.125 200.565 ;
        RECT 32.875 200.020 34.030 200.330 ;
        RECT 32.875 199.745 33.125 200.020 ;
        RECT 11.140 199.575 20.800 199.745 ;
        RECT 23.560 199.575 33.220 199.745 ;
        RECT 36.395 199.725 36.725 200.105 ;
        RECT 37.335 199.725 37.585 200.185 ;
        RECT 39.280 199.725 39.650 200.225 ;
        RECT 41.465 199.725 41.675 200.255 ;
        RECT 42.440 199.725 42.610 200.335 ;
        RECT 43.280 199.725 43.450 200.240 ;
        RECT 44.270 199.725 44.600 200.465 ;
        RECT 45.195 200.380 45.445 200.545 ;
        RECT 45.195 200.010 46.100 200.380 ;
        RECT 135.985 200.090 136.155 201.905 ;
        RECT 45.195 199.725 45.445 200.010 ;
        RECT 35.880 199.555 45.540 199.725 ;
        RECT 135.485 199.720 136.155 200.090 ;
        RECT 135.985 198.025 136.155 199.720 ;
        RECT 135.525 197.775 136.155 198.025 ;
        RECT 135.985 197.165 136.155 197.775 ;
        RECT 135.605 196.835 136.155 197.165 ;
        RECT 135.985 196.320 136.155 196.835 ;
        RECT 96.420 193.870 96.940 194.610 ;
        RECT 97.310 193.870 97.480 194.670 ;
        RECT 96.420 193.825 97.480 193.870 ;
        RECT 98.200 193.825 98.370 194.565 ;
        RECT 99.080 193.825 99.315 194.285 ;
        RECT 101.175 193.825 101.365 194.265 ;
        RECT 103.265 193.825 103.595 194.285 ;
        RECT 106.195 193.825 106.525 194.185 ;
        RECT 107.225 193.825 107.555 194.205 ;
        RECT 96.420 193.655 108.070 193.825 ;
        RECT 96.420 193.640 97.330 193.655 ;
        RECT 136.035 192.635 136.205 192.730 ;
        RECT 135.215 192.385 136.205 192.635 ;
        RECT 136.035 191.790 136.205 192.385 ;
        RECT 135.295 191.460 136.205 191.790 ;
        RECT 136.035 190.640 136.205 191.460 ;
        RECT 135.520 190.470 136.205 190.640 ;
        RECT 98.240 189.480 98.780 190.300 ;
        RECT 98.240 189.475 98.980 189.480 ;
        RECT 100.015 189.475 100.265 189.935 ;
        RECT 101.155 189.475 101.445 190.275 ;
        RECT 98.240 189.305 101.530 189.475 ;
        RECT 103.520 189.455 103.785 189.915 ;
        RECT 104.455 189.455 104.625 189.915 ;
        RECT 105.295 189.455 105.545 189.920 ;
        RECT 136.035 189.800 136.205 190.470 ;
        RECT 135.425 189.630 136.205 189.800 ;
        RECT 98.240 189.300 98.980 189.305 ;
        RECT 103.390 189.285 105.690 189.455 ;
        RECT 136.035 188.865 136.205 189.630 ;
        RECT 135.505 188.655 136.205 188.865 ;
        RECT 136.035 186.840 136.205 188.655 ;
        RECT 135.535 186.470 136.205 186.840 ;
        RECT 96.330 185.090 96.730 185.790 ;
        RECT 97.190 185.090 97.360 185.920 ;
        RECT 96.310 185.075 97.360 185.090 ;
        RECT 98.080 185.075 98.250 185.815 ;
        RECT 98.960 185.075 99.195 185.535 ;
        RECT 101.055 185.075 101.245 185.515 ;
        RECT 103.145 185.075 103.475 185.535 ;
        RECT 106.075 185.075 106.405 185.435 ;
        RECT 107.105 185.075 107.435 185.455 ;
        RECT 96.310 184.905 107.950 185.075 ;
        RECT 96.310 184.900 97.280 184.905 ;
        RECT 136.035 184.775 136.205 186.470 ;
        RECT 135.575 184.525 136.205 184.775 ;
        RECT 136.035 183.915 136.205 184.525 ;
        RECT 135.655 183.585 136.205 183.915 ;
        RECT 136.035 183.210 136.205 183.585 ;
        RECT 136.035 183.070 136.230 183.210 ;
        RECT 136.040 182.900 136.230 183.070 ;
        RECT 135.420 182.380 136.230 182.900 ;
        RECT 121.570 22.190 125.060 22.360 ;
        RECT 121.570 19.090 121.740 22.190 ;
        RECT 121.510 18.320 121.790 19.090 ;
        RECT 121.570 17.540 121.740 18.320 ;
        RECT 122.140 18.220 122.310 21.510 ;
        RECT 124.320 18.220 124.490 21.510 ;
        RECT 124.890 17.540 125.060 22.190 ;
        RECT 140.995 18.225 142.895 18.395 ;
        RECT 121.570 17.370 125.060 17.540 ;
        RECT 137.245 17.765 139.145 17.935 ;
        RECT 99.770 16.820 102.040 16.990 ;
        RECT 99.770 14.440 99.940 16.820 ;
        RECT 99.730 13.920 100.000 14.440 ;
        RECT 99.770 13.170 99.940 13.920 ;
        RECT 100.340 13.850 100.510 16.140 ;
        RECT 101.300 13.850 101.470 16.140 ;
        RECT 101.870 13.170 102.040 16.820 ;
        RECT 104.570 16.890 107.960 17.060 ;
        RECT 104.570 14.600 104.740 16.890 ;
        RECT 104.550 14.010 104.740 14.600 ;
        RECT 99.770 13.000 102.040 13.170 ;
        RECT 104.570 13.240 104.740 14.010 ;
        RECT 107.790 13.240 107.960 16.890 ;
        RECT 104.570 13.070 107.960 13.240 ;
        RECT 110.660 16.870 114.050 17.040 ;
        RECT 110.660 14.530 110.830 16.870 ;
        RECT 110.660 13.970 110.840 14.530 ;
        RECT 110.660 13.220 110.830 13.970 ;
        RECT 113.880 13.220 114.050 16.870 ;
        RECT 116.670 16.880 120.060 17.050 ;
        RECT 116.670 14.470 116.840 16.880 ;
        RECT 116.600 13.970 116.870 14.470 ;
        RECT 110.660 13.050 114.050 13.220 ;
        RECT 116.670 13.230 116.840 13.970 ;
        RECT 119.890 13.230 120.060 16.880 ;
        RECT 137.245 14.365 137.415 17.765 ;
        RECT 138.405 15.045 138.575 17.085 ;
        RECT 138.975 14.365 139.145 17.765 ;
        RECT 140.995 14.840 141.165 18.225 ;
        RECT 142.155 15.505 142.325 17.545 ;
        RECT 140.940 14.825 141.720 14.840 ;
        RECT 142.725 14.825 142.895 18.225 ;
        RECT 140.940 14.655 142.895 14.825 ;
        RECT 144.280 16.260 146.380 16.430 ;
        RECT 140.940 14.400 141.670 14.655 ;
        RECT 137.245 14.360 139.145 14.365 ;
        RECT 137.220 14.195 139.145 14.360 ;
        RECT 140.930 14.340 141.670 14.400 ;
        RECT 141.910 14.340 142.370 14.380 ;
        RECT 137.220 13.980 137.840 14.195 ;
        RECT 140.930 14.070 142.370 14.340 ;
        RECT 144.280 14.200 144.450 16.260 ;
        RECT 145.640 14.840 145.810 15.580 ;
        RECT 144.280 14.160 144.870 14.200 ;
        RECT 146.210 14.160 146.380 16.260 ;
        RECT 137.220 13.820 138.020 13.980 ;
        RECT 140.930 13.970 142.210 14.070 ;
        RECT 144.280 13.990 146.380 14.160 ;
        RECT 140.930 13.960 141.520 13.970 ;
        RECT 137.220 13.640 138.630 13.820 ;
        RECT 144.300 13.740 144.870 13.990 ;
        RECT 116.670 13.060 120.060 13.230 ;
        RECT 137.190 13.200 138.630 13.640 ;
        RECT 138.000 13.100 138.630 13.200 ;
        RECT 143.990 13.180 145.070 13.740 ;
        RECT 148.760 13.290 155.360 13.370 ;
        RECT 145.830 13.200 155.360 13.290 ;
        RECT 145.830 12.770 148.960 13.200 ;
        RECT 146.030 12.690 148.960 12.770 ;
        RECT 104.530 12.030 108.020 12.200 ;
        RECT 104.530 8.950 104.700 12.030 ;
        RECT 104.480 8.110 104.780 8.950 ;
        RECT 104.530 7.380 104.700 8.110 ;
        RECT 105.100 8.060 105.270 11.350 ;
        RECT 107.280 8.060 107.450 11.350 ;
        RECT 107.850 7.380 108.020 12.030 ;
        RECT 110.630 12.030 114.120 12.200 ;
        RECT 110.630 8.970 110.800 12.030 ;
        RECT 110.510 8.130 110.810 8.970 ;
        RECT 104.530 7.210 108.020 7.380 ;
        RECT 110.630 7.380 110.800 8.130 ;
        RECT 111.200 8.060 111.370 11.350 ;
        RECT 113.380 8.060 113.550 11.350 ;
        RECT 113.950 7.380 114.120 12.030 ;
        RECT 116.710 12.050 120.200 12.220 ;
        RECT 116.710 8.820 116.880 12.050 ;
        RECT 116.660 8.170 116.930 8.820 ;
        RECT 110.630 7.210 114.120 7.380 ;
        RECT 116.710 7.400 116.880 8.170 ;
        RECT 117.280 8.080 117.450 11.370 ;
        RECT 119.460 8.080 119.630 11.370 ;
        RECT 120.030 7.400 120.200 12.050 ;
        RECT 148.760 10.800 148.930 12.690 ;
        RECT 155.190 10.800 155.360 13.200 ;
        RECT 148.760 10.630 155.360 10.800 ;
        RECT 116.710 7.230 120.200 7.400 ;
      LAYER met1 ;
        RECT 136.590 220.740 137.590 220.760 ;
        RECT 135.950 219.760 137.590 220.740 ;
        RECT 135.950 219.400 136.320 219.760 ;
        RECT 56.400 217.550 76.840 218.030 ;
        RECT 56.400 214.690 57.060 217.550 ;
        RECT 56.400 214.210 69.020 214.690 ;
        RECT 23.220 214.180 31.960 214.190 ;
        RECT 35.130 214.180 43.870 214.190 ;
        RECT 10.420 214.060 43.870 214.180 ;
        RECT 44.070 214.060 46.460 214.160 ;
        RECT 10.420 213.830 46.460 214.060 ;
        RECT 10.420 213.720 43.870 213.830 ;
        RECT 10.420 213.700 19.160 213.720 ;
        RECT 19.460 213.490 19.760 213.720 ;
        RECT 23.220 213.710 31.960 213.720 ;
        RECT 19.450 213.210 19.770 213.490 ;
        RECT 32.200 213.310 32.620 213.720 ;
        RECT 35.130 213.710 43.870 213.720 ;
        RECT 32.260 213.150 32.580 213.310 ;
        RECT 44.070 212.720 46.460 213.830 ;
        RECT 56.400 211.350 57.060 214.210 ;
        RECT 56.400 210.870 76.840 211.350 ;
        RECT 56.400 202.060 57.400 210.870 ;
        RECT 135.850 209.740 136.330 219.400 ;
        RECT 135.910 205.980 136.190 209.740 ;
        RECT 85.590 202.950 116.330 203.430 ;
        RECT 85.590 202.080 86.590 202.950 ;
        RECT 20.970 200.200 21.430 200.500 ;
        RECT 33.700 200.090 34.040 200.340 ;
        RECT 45.790 199.970 46.110 200.420 ;
        RECT 20.800 199.900 23.680 199.910 ;
        RECT 11.140 199.850 33.220 199.900 ;
        RECT 35.880 199.850 45.540 199.880 ;
        RECT 11.140 199.420 45.540 199.850 ;
        RECT 55.530 199.560 58.130 202.060 ;
        RECT 85.360 199.540 87.220 202.080 ;
        RECT 21.860 199.030 22.990 199.420 ;
        RECT 33.170 199.400 45.540 199.420 ;
        RECT 33.170 199.380 35.970 199.400 ;
        RECT 21.860 198.330 50.440 199.030 ;
        RECT 21.930 198.030 50.440 198.330 ;
        RECT 49.050 196.600 50.350 198.030 ;
        RECT 135.830 196.320 136.310 205.980 ;
        RECT 95.480 193.960 96.490 193.970 ;
        RECT 97.030 193.960 108.070 193.980 ;
        RECT 95.480 193.500 108.070 193.960 ;
        RECT 95.480 189.640 96.490 193.500 ;
        RECT 135.890 192.740 136.310 196.320 ;
        RECT 135.890 192.730 136.370 192.740 ;
        RECT 135.880 192.340 136.370 192.730 ;
        RECT 95.480 189.610 103.770 189.640 ;
        RECT 95.480 189.150 105.690 189.610 ;
        RECT 95.480 185.220 96.490 189.150 ;
        RECT 103.390 189.130 105.690 189.150 ;
        RECT 135.880 186.910 136.360 192.340 ;
        RECT 96.910 185.220 107.950 185.230 ;
        RECT 48.840 184.770 50.740 185.140 ;
        RECT 95.480 184.770 107.950 185.220 ;
        RECT 48.840 184.760 107.950 184.770 ;
        RECT 48.840 183.760 96.515 184.760 ;
        RECT 96.910 184.750 107.950 184.760 ;
        RECT 48.840 183.380 50.740 183.760 ;
        RECT 95.480 183.560 96.490 183.760 ;
        RECT 135.880 183.110 137.940 186.910 ;
        RECT 135.880 183.070 136.360 183.110 ;
        RECT 48.800 180.680 52.490 181.600 ;
        RECT 48.800 180.640 132.650 180.680 ;
        RECT 48.800 180.600 138.010 180.640 ;
        RECT 48.800 178.160 138.040 180.600 ;
        RECT 48.800 177.680 132.650 178.160 ;
        RECT 48.800 177.000 52.490 177.680 ;
        RECT 121.480 19.090 121.820 19.150 ;
        RECT 121.460 18.320 121.840 19.090 ;
        RECT 122.110 19.060 122.340 21.490 ;
        RECT 121.980 18.350 122.430 19.060 ;
        RECT 124.290 19.000 124.520 21.490 ;
        RECT 121.480 18.260 121.820 18.320 ;
        RECT 122.110 18.240 122.340 18.350 ;
        RECT 124.170 18.290 124.620 19.000 ;
        RECT 124.290 18.240 124.520 18.290 ;
        RECT 99.700 14.440 100.030 14.500 ;
        RECT 99.680 13.920 100.050 14.440 ;
        RECT 100.310 14.410 100.540 16.120 ;
        RECT 101.270 14.420 101.500 16.120 ;
        RECT 138.375 15.760 138.605 17.065 ;
        RECT 142.125 16.280 142.355 17.525 ;
        RECT 138.160 15.270 138.790 15.760 ;
        RECT 141.920 15.730 142.660 16.280 ;
        RECT 142.125 15.525 142.355 15.730 ;
        RECT 145.610 15.370 145.840 15.560 ;
        RECT 138.375 15.065 138.605 15.270 ;
        RECT 145.580 14.900 146.270 15.370 ;
        RECT 145.610 14.860 145.840 14.900 ;
        RECT 103.700 14.640 104.120 14.650 ;
        RECT 104.520 14.640 104.770 14.660 ;
        RECT 99.700 13.860 100.030 13.920 ;
        RECT 100.230 13.890 100.600 14.410 ;
        RECT 101.190 13.900 101.560 14.420 ;
        RECT 103.700 13.990 104.840 14.640 ;
        RECT 110.630 14.530 110.870 14.590 ;
        RECT 100.310 13.870 100.540 13.890 ;
        RECT 101.270 13.870 101.500 13.900 ;
        RECT 103.700 12.840 104.120 13.990 ;
        RECT 104.470 13.970 104.840 13.990 ;
        RECT 109.890 14.500 110.370 14.510 ;
        RECT 110.560 14.500 110.940 14.530 ;
        RECT 104.520 13.950 104.770 13.970 ;
        RECT 109.890 13.950 110.940 14.500 ;
        RECT 116.570 14.480 116.900 14.530 ;
        RECT 109.890 12.840 110.370 13.950 ;
        RECT 110.560 13.940 110.940 13.950 ;
        RECT 110.630 13.910 110.870 13.940 ;
        RECT 115.700 13.930 116.920 14.480 ;
        RECT 141.850 14.040 142.430 14.410 ;
        RECT 141.970 14.030 142.350 14.040 ;
        RECT 115.710 12.860 116.350 13.930 ;
        RECT 116.570 13.910 116.900 13.930 ;
        RECT 137.970 13.040 138.660 13.880 ;
        RECT 141.220 13.830 141.670 13.850 ;
        RECT 142.570 13.830 143.090 13.930 ;
        RECT 141.220 13.580 143.090 13.830 ;
        RECT 141.220 13.490 142.780 13.580 ;
        RECT 141.430 13.050 142.780 13.490 ;
        RECT 143.930 13.150 145.130 13.770 ;
        RECT 141.430 12.940 143.090 13.050 ;
        RECT 122.970 12.860 123.600 12.880 ;
        RECT 115.710 12.840 123.600 12.860 ;
        RECT 103.700 12.510 123.600 12.840 ;
        RECT 141.260 12.690 143.090 12.940 ;
        RECT 145.800 12.710 146.350 13.350 ;
        RECT 141.260 12.650 141.700 12.690 ;
        RECT 142.600 12.630 143.090 12.690 ;
        RECT 115.710 12.500 123.600 12.510 ;
        RECT 104.450 8.950 104.810 9.010 ;
        RECT 105.070 8.960 105.300 11.330 ;
        RECT 107.250 8.970 107.480 11.330 ;
        RECT 110.480 8.970 110.840 9.030 ;
        RECT 111.170 9.000 111.400 11.330 ;
        RECT 104.430 8.110 104.830 8.950 ;
        RECT 104.990 8.120 105.390 8.960 ;
        RECT 107.150 8.130 107.550 8.970 ;
        RECT 110.460 8.130 110.860 8.970 ;
        RECT 111.050 8.160 111.450 9.000 ;
        RECT 113.350 8.940 113.580 11.330 ;
        RECT 104.450 8.050 104.810 8.110 ;
        RECT 105.070 8.080 105.300 8.120 ;
        RECT 107.250 8.080 107.480 8.130 ;
        RECT 110.480 8.070 110.840 8.130 ;
        RECT 111.170 8.080 111.400 8.160 ;
        RECT 113.260 8.100 113.660 8.940 ;
        RECT 116.630 8.820 116.960 8.880 ;
        RECT 117.250 8.820 117.480 11.350 ;
        RECT 116.610 8.170 116.980 8.820 ;
        RECT 117.170 8.170 117.540 8.820 ;
        RECT 119.430 8.760 119.660 11.350 ;
        RECT 116.630 8.110 116.960 8.170 ;
        RECT 117.250 8.100 117.480 8.170 ;
        RECT 119.370 8.110 119.740 8.760 ;
        RECT 119.430 8.100 119.660 8.110 ;
        RECT 113.350 8.080 113.580 8.100 ;
        RECT 109.100 6.060 110.210 6.830 ;
        RECT 109.170 5.920 110.170 6.060 ;
        RECT 109.170 4.790 110.430 5.920 ;
        RECT 109.290 3.470 110.430 4.790 ;
        RECT 108.400 2.630 110.960 3.470 ;
      LAYER met2 ;
        RECT 49.000 218.310 50.490 219.000 ;
        RECT 44.120 214.120 46.410 214.210 ;
        RECT 48.910 214.120 50.610 214.420 ;
        RECT 44.120 212.710 50.610 214.120 ;
        RECT 44.120 212.670 46.410 212.710 ;
        RECT 48.910 212.140 50.610 212.710 ;
        RECT 55.580 199.510 58.080 202.110 ;
        RECT 85.410 199.490 87.170 202.130 ;
        RECT 49.100 196.550 50.300 199.010 ;
        RECT 48.890 183.330 50.690 185.190 ;
        RECT 136.200 183.060 137.890 186.960 ;
        RECT 48.850 176.950 52.440 181.650 ;
        RECT 132.650 178.110 137.990 180.650 ;
        RECT 121.510 19.020 121.790 19.140 ;
        RECT 122.030 19.020 122.380 19.110 ;
        RECT 124.220 19.020 124.570 19.050 ;
        RECT 121.500 18.310 124.600 19.020 ;
        RECT 121.510 18.270 121.790 18.310 ;
        RECT 122.030 18.300 122.380 18.310 ;
        RECT 99.730 14.430 100.000 14.490 ;
        RECT 100.280 14.430 100.550 14.460 ;
        RECT 101.240 14.430 101.510 14.470 ;
        RECT 99.700 13.890 101.530 14.430 ;
        RECT 104.520 13.920 104.790 14.690 ;
        RECT 110.610 13.890 110.890 14.580 ;
        RECT 116.600 14.490 116.870 14.520 ;
        RECT 116.540 13.990 116.870 14.490 ;
        RECT 116.600 13.920 116.870 13.990 ;
        RECT 99.730 13.870 100.000 13.890 ;
        RECT 100.280 13.840 100.550 13.890 ;
        RECT 100.750 13.850 101.510 13.890 ;
        RECT 48.970 5.130 52.940 7.460 ;
        RECT 100.750 6.790 101.320 13.850 ;
        RECT 104.480 8.940 104.780 9.000 ;
        RECT 105.040 8.940 105.340 9.010 ;
        RECT 107.200 8.940 107.500 9.020 ;
        RECT 110.510 8.940 110.810 9.020 ;
        RECT 111.100 8.940 111.400 9.050 ;
        RECT 113.310 8.940 113.610 8.990 ;
        RECT 104.420 8.100 119.740 8.940 ;
        RECT 104.480 8.060 104.780 8.100 ;
        RECT 105.040 8.070 105.340 8.100 ;
        RECT 107.200 8.080 107.500 8.100 ;
        RECT 109.140 6.880 110.150 8.100 ;
        RECT 110.510 8.080 110.810 8.100 ;
        RECT 113.310 8.050 113.610 8.100 ;
        RECT 119.420 8.060 119.690 8.100 ;
        RECT 109.140 6.820 110.160 6.880 ;
        RECT 123.010 6.820 123.690 18.310 ;
        RECT 124.220 18.240 124.570 18.310 ;
        RECT 141.970 16.070 142.610 16.330 ;
        RECT 138.190 15.680 138.740 15.810 ;
        RECT 141.970 15.680 142.840 16.070 ;
        RECT 138.190 15.390 139.070 15.680 ;
        RECT 138.190 15.220 139.050 15.390 ;
        RECT 138.340 13.880 139.050 15.220 ;
        RECT 142.110 14.440 142.840 15.680 ;
        RECT 145.630 14.850 146.220 15.420 ;
        RECT 145.630 14.610 146.150 14.850 ;
        RECT 142.020 14.430 142.840 14.440 ;
        RECT 142.020 13.980 142.940 14.430 ;
        RECT 109.140 6.790 123.690 6.820 ;
        RECT 100.750 6.510 123.690 6.790 ;
        RECT 100.780 6.140 123.690 6.510 ;
        RECT 109.150 6.010 123.690 6.140 ;
        RECT 109.430 5.960 123.690 6.010 ;
        RECT 137.940 13.740 139.050 13.880 ;
        RECT 141.270 13.830 141.620 13.900 ;
        RECT 142.110 13.830 143.040 13.980 ;
        RECT 141.270 13.770 143.040 13.830 ;
        RECT 141.270 13.760 143.690 13.770 ;
        RECT 141.270 13.740 143.750 13.760 ;
        RECT 137.940 13.520 143.750 13.740 ;
        RECT 144.200 13.520 144.950 13.720 ;
        RECT 145.600 13.520 146.170 14.610 ;
        RECT 137.940 13.300 146.140 13.520 ;
        RECT 137.940 12.980 146.210 13.300 ;
        RECT 51.660 3.390 52.420 5.130 ;
        RECT 108.450 3.390 110.910 3.520 ;
        RECT 137.940 3.390 138.700 12.980 ;
        RECT 141.270 12.880 146.210 12.980 ;
        RECT 141.270 12.690 143.040 12.880 ;
        RECT 143.600 12.850 143.960 12.880 ;
        RECT 145.930 12.730 146.210 12.880 ;
        RECT 141.270 12.660 141.650 12.690 ;
        RECT 141.310 12.600 141.650 12.660 ;
        RECT 142.650 12.580 143.040 12.690 ;
        RECT 51.660 2.630 138.720 3.390 ;
        RECT 108.450 2.580 110.910 2.630 ;
      LAYER met3 ;
        RECT 22.350 218.790 22.730 218.800 ;
        RECT 48.890 218.790 50.590 219.030 ;
        RECT 22.350 218.490 50.590 218.790 ;
        RECT 22.350 218.480 22.730 218.490 ;
        RECT 48.890 218.280 50.590 218.490 ;
        RECT 48.860 212.165 50.660 214.395 ;
        RECT 48.930 202.060 52.620 202.090 ;
        RECT 55.530 202.060 58.130 202.085 ;
        RECT 85.360 202.060 87.220 202.105 ;
        RECT 48.930 199.560 117.085 202.060 ;
        RECT 55.530 199.535 58.130 199.560 ;
        RECT 85.360 199.515 87.220 199.560 ;
        RECT 49.050 196.575 50.350 198.985 ;
        RECT 136.280 186.935 137.910 186.950 ;
        RECT 48.840 183.355 50.740 185.165 ;
        RECT 136.150 183.085 137.940 186.935 ;
        RECT 48.800 176.975 52.490 181.625 ;
        RECT 136.280 180.625 137.910 183.085 ;
        RECT 132.600 178.135 138.040 180.625 ;
        RECT 48.920 5.155 52.990 7.435 ;
      LAYER met4 ;
        RECT 18.710 218.780 19.010 225.760 ;
        RECT 22.390 218.805 22.690 225.760 ;
        RECT 29.750 220.130 30.050 225.760 ;
        RECT 49.000 220.130 50.500 220.210 ;
        RECT 29.750 219.830 50.500 220.130 ;
        RECT 49.000 219.035 50.500 219.830 ;
        RECT 22.375 218.780 22.705 218.805 ;
        RECT 18.710 218.480 22.810 218.780 ;
        RECT 22.375 218.475 22.705 218.480 ;
        RECT 48.935 218.275 50.545 219.035 ;
        RECT 49.000 214.375 50.500 218.275 ;
        RECT 48.905 212.185 50.615 214.375 ;
        RECT 49.000 202.095 50.500 212.185 ;
        RECT 48.975 199.555 52.575 202.095 ;
        RECT 49.000 185.145 50.500 199.555 ;
        RECT 48.885 183.375 50.695 185.145 ;
        RECT 49.000 181.605 50.500 183.375 ;
        RECT 48.845 176.995 52.445 181.605 ;
        RECT 49.000 7.415 50.500 176.995 ;
        RECT 48.965 5.175 52.945 7.415 ;
        RECT 49.000 5.000 50.500 5.175 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.504000 ;
    ANTENNADIFFAREA 91.085800 ;
    PORT
      LAYER nwell ;
        RECT 56.330 220.700 57.570 220.710 ;
        RECT 56.330 219.260 77.030 220.700 ;
        RECT 57.570 219.095 77.030 219.260 ;
        RECT 133.180 219.590 134.720 220.270 ;
        RECT 62.150 215.910 69.210 217.360 ;
        RECT 63.390 215.755 69.210 215.910 ;
        RECT 10.230 212.580 19.350 212.635 ;
        RECT 10.230 211.510 20.430 212.580 ;
        RECT 23.030 212.540 32.150 212.645 ;
        RECT 10.230 211.030 19.350 211.510 ;
        RECT 23.030 211.500 33.440 212.540 ;
        RECT 34.940 212.000 44.060 212.645 ;
        RECT 59.200 212.570 77.030 214.020 ;
        RECT 60.440 212.415 77.030 212.570 ;
        RECT 23.030 211.040 32.150 211.500 ;
        RECT 34.940 211.040 44.940 212.000 ;
        RECT 43.900 210.890 44.940 211.040 ;
        RECT 133.180 209.550 134.785 219.590 ;
        RECT 85.280 206.100 86.400 206.420 ;
        RECT 133.180 206.170 134.750 209.550 ;
        RECT 85.280 204.890 116.520 206.100 ;
        RECT 86.400 204.495 116.520 204.890 ;
        RECT 10.950 201.730 21.590 202.570 ;
        RECT 23.370 202.560 33.410 202.570 ;
        RECT 10.950 200.965 20.990 201.730 ;
        RECT 23.370 201.220 34.370 202.560 ;
        RECT 45.720 202.550 47.100 202.560 ;
        RECT 23.370 200.965 33.410 201.220 ;
        RECT 35.690 200.960 47.100 202.550 ;
        RECT 35.690 200.945 45.730 200.960 ;
        RECT 95.710 196.650 97.250 196.690 ;
        RECT 95.710 195.045 108.260 196.650 ;
        RECT 133.160 196.290 134.765 206.170 ;
        RECT 133.160 196.130 134.790 196.290 ;
        RECT 95.710 195.000 97.250 195.045 ;
        RECT 133.200 192.920 134.790 196.130 ;
        RECT 133.200 192.740 134.815 192.920 ;
        RECT 97.860 192.300 98.770 192.310 ;
        RECT 97.860 192.280 103.320 192.300 ;
        RECT 97.860 191.320 105.880 192.280 ;
        RECT 98.580 190.695 105.880 191.320 ;
        RECT 101.540 190.680 105.880 190.695 ;
        RECT 103.200 190.675 105.880 190.680 ;
        RECT 95.930 187.900 97.020 187.970 ;
        RECT 95.930 186.295 108.140 187.900 ;
        RECT 95.930 186.240 97.020 186.295 ;
        RECT 133.210 182.880 134.815 192.740 ;
        RECT 106.070 23.170 109.920 28.610 ;
        RECT 111.190 23.170 115.040 28.610 ;
        RECT 116.310 23.160 120.160 28.600 ;
        RECT 121.430 23.160 125.280 28.600 ;
        RECT 99.220 17.770 102.330 21.960 ;
        RECT 103.610 17.710 108.400 21.900 ;
        RECT 109.670 17.710 114.460 21.900 ;
        RECT 115.730 17.700 120.520 21.890 ;
        RECT 138.850 19.580 142.290 27.770 ;
        RECT 144.600 19.260 146.860 27.450 ;
        RECT 150.880 18.810 153.730 28.000 ;
        RECT 150.285 14.340 154.245 17.530 ;
      LAYER li1 ;
        RECT 56.560 220.595 57.760 220.630 ;
        RECT 56.560 220.425 60.060 220.595 ;
        RECT 60.440 220.425 62.740 220.595 ;
        RECT 63.120 220.425 65.420 220.595 ;
        RECT 65.800 220.425 76.840 220.595 ;
        RECT 56.560 220.420 57.760 220.425 ;
        RECT 56.560 219.510 57.390 220.420 ;
        RECT 57.945 219.965 58.155 220.425 ;
        RECT 58.825 219.625 58.995 220.425 ;
        RECT 59.665 219.285 59.930 220.425 ;
        RECT 60.625 219.965 60.835 220.425 ;
        RECT 61.505 219.625 61.675 220.425 ;
        RECT 62.345 219.285 62.610 220.425 ;
        RECT 63.305 219.965 63.515 220.425 ;
        RECT 64.185 219.625 64.355 220.425 ;
        RECT 65.025 219.285 65.290 220.425 ;
        RECT 66.080 219.235 66.250 220.425 ;
        RECT 66.890 220.045 67.220 220.425 ;
        RECT 67.770 219.995 68.110 220.425 ;
        RECT 68.785 220.045 69.130 220.425 ;
        RECT 69.650 219.965 69.900 220.425 ;
        RECT 71.515 219.965 71.885 220.425 ;
        RECT 72.520 219.995 72.850 220.425 ;
        RECT 74.740 219.965 74.990 220.425 ;
        RECT 75.240 220.240 75.430 220.425 ;
        RECT 75.160 219.455 75.485 220.240 ;
        RECT 75.995 219.925 76.325 220.425 ;
        RECT 133.250 220.080 134.540 220.110 ;
        RECT 133.210 219.580 134.540 220.080 ;
        RECT 74.965 218.405 75.425 219.455 ;
        RECT 133.210 219.350 133.490 219.580 ;
        RECT 133.280 219.305 133.490 219.350 ;
        RECT 133.280 219.250 134.595 219.305 ;
        RECT 133.285 219.055 134.595 219.250 ;
        RECT 133.285 218.380 133.455 219.055 ;
        RECT 133.285 218.165 134.595 218.380 ;
        RECT 133.285 217.305 133.455 218.165 ;
        RECT 62.380 217.255 63.580 217.280 ;
        RECT 62.380 217.085 66.340 217.255 ;
        RECT 66.720 217.085 69.020 217.255 ;
        RECT 133.285 217.130 134.370 217.305 ;
        RECT 62.380 217.080 63.580 217.085 ;
        RECT 62.380 216.160 63.210 217.080 ;
        RECT 63.865 216.415 64.145 217.085 ;
        RECT 64.825 216.365 65.155 217.085 ;
        RECT 65.965 215.945 66.255 217.085 ;
        RECT 66.850 215.945 67.115 217.085 ;
        RECT 67.785 216.285 67.955 217.085 ;
        RECT 68.625 216.625 68.835 217.085 ;
        RECT 133.285 216.460 133.455 217.130 ;
        RECT 133.285 216.290 134.465 216.460 ;
        RECT 133.285 215.545 133.455 216.290 ;
        RECT 133.285 215.230 133.955 215.545 ;
        RECT 59.430 213.915 60.630 213.930 ;
        RECT 59.430 213.745 62.930 213.915 ;
        RECT 63.310 213.745 65.610 213.915 ;
        RECT 65.800 213.745 76.840 213.915 ;
        RECT 59.430 213.740 60.630 213.745 ;
        RECT 59.430 212.820 60.260 213.740 ;
        RECT 60.815 213.285 61.025 213.745 ;
        RECT 61.695 212.945 61.865 213.745 ;
        RECT 62.535 212.605 62.800 213.745 ;
        RECT 63.495 213.285 63.705 213.745 ;
        RECT 64.375 212.945 64.545 213.745 ;
        RECT 65.215 212.605 65.480 213.745 ;
        RECT 66.080 212.555 66.250 213.745 ;
        RECT 66.890 213.365 67.220 213.745 ;
        RECT 67.770 213.315 68.110 213.745 ;
        RECT 68.785 213.365 69.130 213.745 ;
        RECT 69.650 213.285 69.900 213.745 ;
        RECT 71.515 213.285 71.885 213.745 ;
        RECT 72.520 213.315 72.850 213.745 ;
        RECT 74.740 213.285 74.990 213.745 ;
        RECT 75.230 213.560 75.420 213.745 ;
        RECT 75.160 212.775 75.485 213.560 ;
        RECT 75.995 213.245 76.325 213.745 ;
        RECT 133.285 213.520 133.455 215.230 ;
        RECT 133.285 213.350 134.255 213.520 ;
        RECT 10.935 211.305 11.265 211.805 ;
        RECT 11.860 211.305 12.125 211.765 ;
        RECT 14.030 211.305 14.200 212.105 ;
        RECT 15.910 211.305 16.225 211.805 ;
        RECT 16.970 211.305 17.140 212.315 ;
        RECT 18.350 211.305 18.565 212.445 ;
        RECT 19.370 211.740 19.800 212.360 ;
        RECT 10.420 211.300 19.160 211.305 ;
        RECT 19.460 211.300 19.650 211.740 ;
        RECT 23.735 211.315 24.065 211.815 ;
        RECT 24.660 211.315 24.925 211.775 ;
        RECT 26.830 211.315 27.000 212.115 ;
        RECT 28.710 211.315 29.025 211.815 ;
        RECT 29.770 211.315 29.940 212.325 ;
        RECT 31.150 211.315 31.365 212.455 ;
        RECT 32.170 211.720 32.640 212.280 ;
        RECT 10.420 211.135 19.650 211.300 ;
        RECT 23.220 211.310 31.960 211.315 ;
        RECT 32.200 211.310 32.420 211.720 ;
        RECT 35.645 211.315 35.975 211.815 ;
        RECT 36.570 211.315 36.835 211.775 ;
        RECT 38.740 211.315 38.910 212.115 ;
        RECT 40.620 211.315 40.935 211.815 ;
        RECT 41.680 211.315 41.850 212.325 ;
        RECT 43.060 211.315 43.275 212.455 ;
        RECT 23.220 211.145 32.420 211.310 ;
        RECT 35.130 211.310 43.870 211.315 ;
        RECT 44.180 211.310 44.450 211.780 ;
        RECT 74.965 211.725 75.425 212.775 ;
        RECT 35.130 211.145 44.450 211.310 ;
        RECT 31.650 211.140 32.420 211.145 ;
        RECT 43.550 211.140 44.450 211.145 ;
        RECT 18.810 211.110 19.650 211.135 ;
        RECT 32.200 211.130 32.420 211.140 ;
        RECT 44.180 211.120 44.450 211.140 ;
        RECT 133.285 211.445 133.455 213.350 ;
        RECT 133.285 211.180 133.915 211.445 ;
        RECT 133.285 210.585 133.455 211.180 ;
        RECT 133.285 210.255 133.955 210.585 ;
        RECT 133.285 209.740 133.455 210.255 ;
        RECT 85.640 206.020 86.150 206.180 ;
        RECT 85.640 205.830 87.970 206.020 ;
        RECT 85.640 205.140 86.150 205.830 ;
        RECT 86.590 205.825 87.970 205.830 ;
        RECT 88.160 205.825 89.540 205.995 ;
        RECT 89.770 205.825 98.510 205.995 ;
        RECT 98.680 205.825 107.420 205.995 ;
        RECT 107.590 205.825 116.330 205.995 ;
        RECT 133.265 205.885 133.435 205.980 ;
        RECT 86.735 204.685 86.945 205.825 ;
        RECT 87.615 204.685 87.845 205.825 ;
        RECT 88.305 204.685 88.515 205.825 ;
        RECT 89.185 204.685 89.415 205.825 ;
        RECT 90.365 204.685 90.580 205.825 ;
        RECT 91.790 204.815 91.960 205.825 ;
        RECT 92.705 205.325 93.020 205.825 ;
        RECT 94.730 205.025 94.900 205.825 ;
        RECT 96.805 205.365 97.070 205.825 ;
        RECT 97.665 205.325 97.995 205.825 ;
        RECT 99.275 204.685 99.490 205.825 ;
        RECT 100.700 204.815 100.870 205.825 ;
        RECT 101.615 205.325 101.930 205.825 ;
        RECT 103.640 205.025 103.810 205.825 ;
        RECT 105.715 205.365 105.980 205.825 ;
        RECT 106.575 205.325 106.905 205.825 ;
        RECT 108.185 204.685 108.400 205.825 ;
        RECT 109.610 204.815 109.780 205.825 ;
        RECT 110.525 205.325 110.840 205.825 ;
        RECT 112.550 205.025 112.720 205.825 ;
        RECT 114.625 205.365 114.890 205.825 ;
        RECT 115.485 205.325 115.815 205.825 ;
        RECT 133.265 205.635 134.575 205.885 ;
        RECT 133.265 204.960 133.435 205.635 ;
        RECT 133.265 204.745 134.575 204.960 ;
        RECT 133.265 203.885 133.435 204.745 ;
        RECT 133.265 203.710 134.350 203.885 ;
        RECT 133.265 203.040 133.435 203.710 ;
        RECT 133.265 202.870 134.445 203.040 ;
        RECT 20.480 202.465 20.800 202.470 ;
        RECT 11.140 202.295 20.800 202.465 ;
        RECT 23.560 202.295 33.220 202.465 ;
        RECT 11.655 201.795 11.985 202.295 ;
        RECT 12.580 201.835 12.845 202.295 ;
        RECT 14.750 201.495 14.920 202.295 ;
        RECT 16.630 201.795 16.945 202.295 ;
        RECT 17.690 201.285 17.860 202.295 ;
        RECT 18.530 201.380 18.705 202.295 ;
        RECT 19.565 201.155 19.780 202.295 ;
        RECT 20.455 202.260 20.800 202.295 ;
        RECT 20.455 202.000 21.360 202.260 ;
        RECT 20.455 201.155 20.705 202.000 ;
        RECT 24.075 201.795 24.405 202.295 ;
        RECT 25.000 201.835 25.265 202.295 ;
        RECT 27.170 201.495 27.340 202.295 ;
        RECT 29.050 201.795 29.365 202.295 ;
        RECT 30.110 201.285 30.280 202.295 ;
        RECT 30.950 201.380 31.125 202.295 ;
        RECT 31.985 201.155 32.200 202.295 ;
        RECT 32.875 201.990 33.125 202.295 ;
        RECT 35.880 202.275 45.540 202.445 ;
        RECT 32.875 201.650 34.030 201.990 ;
        RECT 36.395 201.775 36.725 202.275 ;
        RECT 37.320 201.815 37.585 202.275 ;
        RECT 32.875 201.155 33.125 201.650 ;
        RECT 39.490 201.475 39.660 202.275 ;
        RECT 41.370 201.775 41.685 202.275 ;
        RECT 42.430 201.265 42.600 202.275 ;
        RECT 43.270 201.360 43.445 202.275 ;
        RECT 44.305 201.135 44.520 202.275 ;
        RECT 45.195 202.010 45.445 202.275 ;
        RECT 133.265 202.125 133.435 202.870 ;
        RECT 45.195 201.570 46.690 202.010 ;
        RECT 133.265 201.810 133.935 202.125 ;
        RECT 45.195 201.135 45.445 201.570 ;
        RECT 133.265 200.100 133.435 201.810 ;
        RECT 133.265 199.930 134.235 200.100 ;
        RECT 133.265 198.025 133.435 199.930 ;
        RECT 133.265 197.760 133.895 198.025 ;
        RECT 133.265 197.165 133.435 197.760 ;
        RECT 133.265 196.835 133.935 197.165 ;
        RECT 96.530 196.550 96.880 196.570 ;
        RECT 96.530 196.545 97.090 196.550 ;
        RECT 96.530 196.375 108.070 196.545 ;
        RECT 96.530 196.370 97.090 196.375 ;
        RECT 96.530 195.600 96.880 196.370 ;
        RECT 97.310 195.185 97.480 196.375 ;
        RECT 98.120 195.995 98.450 196.375 ;
        RECT 99.000 195.945 99.340 196.375 ;
        RECT 100.015 195.995 100.360 196.375 ;
        RECT 100.880 195.915 101.130 196.375 ;
        RECT 102.745 195.915 103.115 196.375 ;
        RECT 103.750 195.945 104.080 196.375 ;
        RECT 105.970 195.915 106.220 196.375 ;
        RECT 106.420 196.190 106.680 196.375 ;
        RECT 106.390 195.405 106.715 196.190 ;
        RECT 107.225 195.875 107.555 196.375 ;
        RECT 133.265 196.320 133.435 196.835 ;
        RECT 106.195 194.355 106.655 195.405 ;
        RECT 133.315 192.635 133.485 192.730 ;
        RECT 133.315 192.385 134.625 192.635 ;
        RECT 98.070 192.195 98.830 192.220 ;
        RECT 98.070 192.025 101.530 192.195 ;
        RECT 98.070 192.000 98.830 192.025 ;
        RECT 98.070 191.550 98.440 192.000 ;
        RECT 99.055 191.355 99.335 192.025 ;
        RECT 100.015 191.305 100.345 192.025 ;
        RECT 101.155 190.885 101.445 192.025 ;
        RECT 103.390 192.005 105.690 192.175 ;
        RECT 103.520 190.865 103.785 192.005 ;
        RECT 104.455 191.205 104.625 192.005 ;
        RECT 105.295 191.545 105.505 192.005 ;
        RECT 133.315 191.710 133.485 192.385 ;
        RECT 133.315 191.495 134.625 191.710 ;
        RECT 133.315 190.635 133.485 191.495 ;
        RECT 133.315 190.460 134.400 190.635 ;
        RECT 133.315 189.790 133.485 190.460 ;
        RECT 133.315 189.620 134.495 189.790 ;
        RECT 133.315 188.875 133.485 189.620 ;
        RECT 133.315 188.560 133.985 188.875 ;
        RECT 96.270 187.795 96.990 187.820 ;
        RECT 96.270 187.625 107.950 187.795 ;
        RECT 96.270 187.590 96.990 187.625 ;
        RECT 96.290 186.710 96.700 187.590 ;
        RECT 97.190 186.435 97.360 187.625 ;
        RECT 98.000 187.245 98.330 187.625 ;
        RECT 98.880 187.195 99.220 187.625 ;
        RECT 99.895 187.245 100.240 187.625 ;
        RECT 100.760 187.165 101.010 187.625 ;
        RECT 102.625 187.165 102.995 187.625 ;
        RECT 103.630 187.195 103.960 187.625 ;
        RECT 105.850 187.165 106.100 187.625 ;
        RECT 106.310 187.440 106.570 187.625 ;
        RECT 106.270 186.655 106.595 187.440 ;
        RECT 107.105 187.125 107.435 187.625 ;
        RECT 133.315 186.850 133.485 188.560 ;
        RECT 133.315 186.680 134.285 186.850 ;
        RECT 106.075 185.605 106.535 186.655 ;
        RECT 133.315 184.775 133.485 186.680 ;
        RECT 133.315 184.510 133.945 184.775 ;
        RECT 133.315 183.915 133.485 184.510 ;
        RECT 133.315 183.585 133.985 183.915 ;
        RECT 133.315 183.070 133.485 183.585 ;
        RECT 151.870 29.320 152.970 29.530 ;
        RECT 106.250 28.260 109.740 28.430 ;
        RECT 106.250 27.510 106.420 28.260 ;
        RECT 106.220 26.860 106.510 27.510 ;
        RECT 106.250 23.520 106.420 26.860 ;
        RECT 106.820 24.245 106.990 27.535 ;
        RECT 109.000 24.245 109.170 27.535 ;
        RECT 109.570 23.520 109.740 28.260 ;
        RECT 111.370 28.260 114.860 28.430 ;
        RECT 111.370 27.400 111.540 28.260 ;
        RECT 111.320 26.700 111.610 27.400 ;
        RECT 106.250 23.350 109.740 23.520 ;
        RECT 111.370 23.520 111.540 26.700 ;
        RECT 111.940 24.245 112.110 27.535 ;
        RECT 114.120 24.245 114.290 27.535 ;
        RECT 114.690 23.520 114.860 28.260 ;
        RECT 116.490 28.250 119.980 28.420 ;
        RECT 116.490 27.390 116.660 28.250 ;
        RECT 116.480 26.770 116.670 27.390 ;
        RECT 111.370 23.350 114.860 23.520 ;
        RECT 116.490 23.510 116.660 26.770 ;
        RECT 117.060 24.235 117.230 27.525 ;
        RECT 119.240 24.235 119.410 27.525 ;
        RECT 119.810 23.510 119.980 28.250 ;
        RECT 121.610 28.250 125.100 28.420 ;
        RECT 121.610 27.470 121.780 28.250 ;
        RECT 121.570 26.820 121.800 27.470 ;
        RECT 116.490 23.340 119.980 23.510 ;
        RECT 121.610 23.510 121.780 26.820 ;
        RECT 122.180 24.235 122.350 27.525 ;
        RECT 124.360 24.235 124.530 27.525 ;
        RECT 124.930 23.510 125.100 28.250 ;
        RECT 143.230 27.820 145.210 28.410 ;
        RECT 151.870 28.090 153.640 29.320 ;
        RECT 152.970 27.820 153.640 28.090 ;
        RECT 121.610 23.340 125.100 23.510 ;
        RECT 139.030 27.580 142.110 27.590 ;
        RECT 143.700 27.580 144.950 27.820 ;
        RECT 139.030 27.420 144.950 27.580 ;
        RECT 99.400 21.610 102.150 21.780 ;
        RECT 99.400 20.860 99.570 21.610 ;
        RECT 99.300 20.430 99.620 20.860 ;
        RECT 99.400 18.120 99.570 20.430 ;
        RECT 100.450 18.845 100.620 20.885 ;
        RECT 101.410 18.845 101.580 20.885 ;
        RECT 101.980 18.120 102.150 21.610 ;
        RECT 103.790 21.550 108.220 21.720 ;
        RECT 103.790 20.830 103.960 21.550 ;
        RECT 103.780 20.400 103.980 20.830 ;
        RECT 99.400 17.950 102.150 18.120 ;
        RECT 103.790 18.060 103.960 20.400 ;
        RECT 108.050 18.060 108.220 21.550 ;
        RECT 109.850 21.550 114.280 21.720 ;
        RECT 109.850 20.790 110.020 21.550 ;
        RECT 109.810 20.380 110.080 20.790 ;
        RECT 103.790 17.890 108.220 18.060 ;
        RECT 109.850 18.060 110.020 20.380 ;
        RECT 114.110 18.060 114.280 21.550 ;
        RECT 115.910 21.540 120.340 21.710 ;
        RECT 115.910 20.770 116.080 21.540 ;
        RECT 115.850 20.230 116.110 20.770 ;
        RECT 109.850 17.890 114.280 18.060 ;
        RECT 115.910 18.050 116.080 20.230 ;
        RECT 120.170 18.050 120.340 21.540 ;
        RECT 139.030 19.930 139.200 27.420 ;
        RECT 141.830 27.270 144.950 27.420 ;
        RECT 151.060 27.650 153.640 27.820 ;
        RECT 141.830 27.100 146.680 27.270 ;
        RECT 141.830 26.790 144.950 27.100 ;
        RECT 140.190 20.655 140.360 26.695 ;
        RECT 141.370 20.655 141.540 26.695 ;
        RECT 141.830 26.220 144.970 26.790 ;
        RECT 141.940 19.930 142.110 26.220 ;
        RECT 143.710 26.180 144.970 26.220 ;
        RECT 139.030 19.760 142.110 19.930 ;
        RECT 144.780 19.610 144.950 26.180 ;
        RECT 145.940 20.335 146.110 26.375 ;
        RECT 146.510 19.610 146.680 27.100 ;
        RECT 144.780 19.440 146.680 19.610 ;
        RECT 151.060 19.160 151.230 27.650 ;
        RECT 152.970 27.170 153.640 27.650 ;
        RECT 152.220 19.885 152.390 26.925 ;
        RECT 153.380 19.160 153.550 27.170 ;
        RECT 151.060 18.990 153.550 19.160 ;
        RECT 115.910 17.880 120.340 18.050 ;
        RECT 151.080 17.350 152.130 18.990 ;
        RECT 150.465 17.180 154.065 17.350 ;
        RECT 150.465 14.690 150.635 17.180 ;
        RECT 153.895 14.690 154.065 17.180 ;
        RECT 150.465 14.520 154.065 14.690 ;
      LAYER met1 ;
        RECT 77.370 220.750 78.370 221.750 ;
        RECT 57.410 220.280 78.370 220.750 ;
        RECT 57.410 220.270 65.420 220.280 ;
        RECT 65.800 220.270 78.370 220.280 ;
        RECT 77.710 217.650 78.370 220.270 ;
        RECT 77.620 217.410 78.430 217.650 ;
        RECT 63.580 216.930 78.430 217.410 ;
        RECT 77.620 214.070 78.430 216.930 ;
        RECT 59.670 213.760 78.430 214.070 ;
        RECT 59.670 213.600 78.370 213.760 ;
        RECT 60.630 213.590 62.930 213.600 ;
        RECT 63.310 213.590 65.610 213.600 ;
        RECT 65.800 213.590 78.370 213.600 ;
        RECT 9.120 211.010 43.870 211.470 ;
        RECT 9.140 210.980 19.160 211.010 ;
        RECT 23.220 210.990 31.960 211.010 ;
        RECT 35.130 210.990 43.870 211.010 ;
        RECT 9.140 209.060 11.990 210.980 ;
        RECT 133.130 209.740 133.610 219.400 ;
        RECT 9.070 206.560 12.260 209.060 ;
        RECT 21.960 208.790 22.960 208.820 ;
        RECT 19.220 206.880 25.350 208.790 ;
        RECT 21.960 203.540 22.960 206.880 ;
        RECT 82.120 206.660 84.040 209.000 ;
        RECT 21.950 203.120 22.960 203.540 ;
        RECT 21.950 202.620 22.950 203.120 ;
        RECT 11.130 202.600 36.020 202.620 ;
        RECT 11.130 202.150 45.540 202.600 ;
        RECT 11.130 202.140 33.220 202.150 ;
        RECT 11.130 202.120 33.190 202.140 ;
        RECT 35.880 202.120 45.540 202.150 ;
        RECT 82.460 198.200 83.460 206.660 ;
        RECT 114.990 206.150 117.360 209.140 ;
        RECT 86.590 205.670 117.360 206.150 ;
        RECT 133.210 205.980 133.490 209.740 ;
        RECT 82.460 197.200 109.410 198.200 ;
        RECT 108.340 196.700 109.340 197.200 ;
        RECT 97.030 196.240 109.340 196.700 ;
        RECT 133.110 196.320 133.590 205.980 ;
        RECT 97.030 196.220 108.070 196.240 ;
        RECT 98.770 192.340 101.530 192.350 ;
        RECT 98.770 192.330 103.710 192.340 ;
        RECT 105.200 192.330 105.740 192.340 ;
        RECT 98.770 191.890 105.740 192.330 ;
        RECT 98.770 191.870 101.530 191.890 ;
        RECT 103.390 191.880 105.740 191.890 ;
        RECT 103.390 191.850 105.690 191.880 ;
        RECT 96.910 187.940 107.950 187.950 ;
        RECT 108.290 187.940 109.340 196.240 ;
        RECT 133.170 192.730 133.590 196.320 ;
        RECT 96.910 187.480 109.340 187.940 ;
        RECT 96.910 187.470 107.950 187.480 ;
        RECT 133.160 183.480 133.640 192.730 ;
        RECT 133.150 183.070 133.640 183.480 ;
        RECT 125.070 182.430 129.510 182.500 ;
        RECT 133.150 182.430 133.620 183.070 ;
        RECT 125.070 181.430 133.620 182.430 ;
        RECT 125.070 181.410 129.510 181.430 ;
        RECT 113.050 31.700 118.240 33.150 ;
        RECT 115.030 30.520 116.420 31.700 ;
        RECT 114.920 29.630 116.420 30.520 ;
        RECT 114.920 29.520 115.920 29.630 ;
        RECT 115.060 29.380 115.840 29.520 ;
        RECT 115.030 28.640 115.880 29.380 ;
        RECT 144.440 28.660 145.740 29.890 ;
        RECT 143.170 27.790 145.270 28.440 ;
        RECT 151.840 28.030 153.000 29.590 ;
        RECT 106.190 27.510 106.540 27.570 ;
        RECT 106.170 26.860 106.560 27.510 ;
        RECT 106.790 27.450 107.020 27.515 ;
        RECT 108.970 27.470 109.200 27.515 ;
        RECT 111.910 27.480 112.140 27.515 ;
        RECT 106.190 26.800 106.540 26.860 ;
        RECT 106.740 26.820 107.100 27.450 ;
        RECT 108.960 26.840 109.320 27.470 ;
        RECT 111.290 27.400 111.640 27.460 ;
        RECT 106.790 24.265 107.020 26.820 ;
        RECT 108.970 24.265 109.200 26.840 ;
        RECT 111.270 26.700 111.660 27.400 ;
        RECT 111.800 26.780 112.190 27.480 ;
        RECT 114.090 27.440 114.320 27.515 ;
        RECT 111.290 26.640 111.640 26.700 ;
        RECT 111.910 24.265 112.140 26.780 ;
        RECT 114.060 26.740 114.450 27.440 ;
        RECT 114.090 24.265 114.320 26.740 ;
        RECT 116.350 26.710 116.750 27.500 ;
        RECT 117.030 27.480 117.260 27.505 ;
        RECT 116.950 26.850 117.310 27.480 ;
        RECT 119.210 27.440 119.440 27.505 ;
        RECT 117.030 24.255 117.260 26.850 ;
        RECT 119.140 26.810 119.500 27.440 ;
        RECT 119.210 24.255 119.440 26.810 ;
        RECT 121.480 26.760 121.890 27.530 ;
        RECT 122.090 26.880 122.450 27.510 ;
        RECT 124.280 26.880 124.640 27.510 ;
        RECT 122.150 24.255 122.380 26.880 ;
        RECT 124.330 24.255 124.560 26.880 ;
        RECT 140.160 26.320 140.390 26.675 ;
        RECT 140.030 25.040 140.530 26.320 ;
        RECT 141.340 26.310 141.570 26.675 ;
        RECT 152.190 26.420 152.420 26.905 ;
        RECT 103.680 23.060 104.190 23.150 ;
        RECT 109.660 23.060 110.190 23.070 ;
        RECT 103.680 22.760 116.270 23.060 ;
        RECT 103.830 22.740 116.270 22.760 ;
        RECT 99.270 20.860 99.650 20.920 ;
        RECT 100.420 20.860 100.650 20.865 ;
        RECT 99.250 20.430 99.670 20.860 ;
        RECT 100.330 20.430 100.750 20.860 ;
        RECT 101.280 20.440 101.700 20.870 ;
        RECT 103.750 20.840 104.010 20.890 ;
        RECT 99.270 20.370 99.650 20.430 ;
        RECT 100.420 18.865 100.650 20.430 ;
        RECT 101.380 18.865 101.610 20.440 ;
        RECT 103.690 20.370 104.050 20.840 ;
        RECT 109.780 20.790 110.110 20.850 ;
        RECT 109.760 20.380 110.130 20.790 ;
        RECT 115.820 20.770 116.140 20.830 ;
        RECT 103.750 20.340 104.010 20.370 ;
        RECT 109.780 20.320 110.110 20.380 ;
        RECT 115.800 20.230 116.160 20.770 ;
        RECT 140.160 20.675 140.390 25.040 ;
        RECT 141.190 25.030 141.690 26.310 ;
        RECT 145.910 26.130 146.140 26.355 ;
        RECT 145.790 25.520 146.330 26.130 ;
        RECT 141.340 20.675 141.570 25.030 ;
        RECT 145.910 20.355 146.140 25.520 ;
        RECT 152.110 25.320 152.550 26.420 ;
        RECT 115.820 20.170 116.140 20.230 ;
        RECT 152.190 19.905 152.420 25.320 ;
      LAYER met2 ;
        RECT 77.670 213.710 78.380 217.700 ;
        RECT 9.120 206.510 12.210 209.110 ;
        RECT 19.270 206.830 25.300 208.840 ;
        RECT 82.170 206.610 83.990 209.050 ;
        RECT 115.040 205.620 117.310 209.190 ;
        RECT 105.250 192.340 105.690 192.390 ;
        RECT 108.700 192.340 109.140 192.370 ;
        RECT 105.250 191.860 109.140 192.340 ;
        RECT 105.250 191.830 105.690 191.860 ;
        RECT 108.700 191.810 109.140 191.860 ;
        RECT 125.120 181.360 129.460 182.550 ;
        RECT 1.010 32.995 5.080 33.890 ;
        RECT 113.100 32.995 118.190 33.200 ;
        RECT 1.010 32.980 142.075 32.995 ;
        RECT 1.010 31.725 142.130 32.980 ;
        RECT 1.010 30.360 5.080 31.725 ;
        RECT 113.100 31.650 118.190 31.725 ;
        RECT 100.630 29.460 101.350 29.480 ;
        RECT 100.630 29.430 115.740 29.460 ;
        RECT 100.630 29.060 115.830 29.430 ;
        RECT 140.180 29.300 142.130 31.725 ;
        RECT 144.130 29.300 145.850 29.960 ;
        RECT 152.020 29.330 152.820 29.460 ;
        RECT 147.550 29.300 152.820 29.330 ;
        RECT 100.630 28.700 115.840 29.060 ;
        RECT 100.630 20.920 101.350 28.700 ;
        RECT 103.680 22.760 104.140 28.700 ;
        RECT 106.220 27.510 106.510 27.560 ;
        RECT 109.010 27.510 109.270 27.520 ;
        RECT 111.850 27.510 112.140 27.530 ;
        RECT 115.080 27.510 115.840 28.700 ;
        RECT 140.180 28.060 152.820 29.300 ;
        RECT 140.550 28.040 152.770 28.060 ;
        RECT 116.400 27.510 116.700 27.550 ;
        RECT 117.000 27.510 117.260 27.530 ;
        RECT 121.530 27.510 121.840 27.580 ;
        RECT 122.140 27.510 122.400 27.560 ;
        RECT 124.330 27.510 124.590 27.560 ;
        RECT 106.220 26.880 124.680 27.510 ;
        RECT 106.220 26.810 106.510 26.880 ;
        RECT 106.790 26.770 107.050 26.880 ;
        RECT 109.010 26.790 109.270 26.880 ;
        RECT 111.320 26.650 111.610 26.880 ;
        RECT 111.850 26.730 112.140 26.880 ;
        RECT 114.110 26.690 114.400 26.880 ;
        RECT 116.400 26.660 116.700 26.880 ;
        RECT 117.000 26.800 117.260 26.880 ;
        RECT 119.190 26.760 119.450 26.880 ;
        RECT 121.530 26.710 121.840 26.880 ;
        RECT 122.140 26.830 122.400 26.880 ;
        RECT 124.330 26.830 124.590 26.880 ;
        RECT 140.550 26.570 141.760 28.040 ;
        RECT 143.470 27.870 145.130 28.040 ;
        RECT 140.390 26.370 141.760 26.570 ;
        RECT 140.080 26.270 141.760 26.370 ;
        RECT 139.910 25.080 141.760 26.270 ;
        RECT 145.890 26.180 146.760 28.040 ;
        RECT 147.550 28.030 152.770 28.040 ;
        RECT 151.750 27.310 152.770 28.030 ;
        RECT 151.750 27.300 152.780 27.310 ;
        RECT 145.840 25.670 146.760 26.180 ;
        RECT 151.780 26.430 152.780 27.300 ;
        RECT 145.840 25.470 146.280 25.670 ;
        RECT 151.780 25.320 152.820 26.430 ;
        RECT 152.160 25.270 152.500 25.320 ;
        RECT 140.080 25.020 141.760 25.080 ;
        RECT 140.080 24.990 140.670 25.020 ;
        RECT 140.410 24.970 140.670 24.990 ;
        RECT 141.240 24.980 141.640 25.020 ;
        RECT 103.720 22.710 104.140 22.760 ;
        RECT 100.630 20.910 101.650 20.920 ;
        RECT 99.300 20.870 99.620 20.910 ;
        RECT 100.380 20.870 101.650 20.910 ;
        RECT 99.290 20.440 101.710 20.870 ;
        RECT 99.300 20.380 99.620 20.440 ;
        RECT 100.380 20.380 100.700 20.440 ;
        RECT 101.330 20.390 101.650 20.440 ;
        RECT 103.720 20.390 104.110 22.710 ;
        RECT 109.710 22.700 110.140 23.120 ;
        RECT 103.740 20.320 104.000 20.390 ;
        RECT 109.740 20.330 110.130 22.700 ;
        RECT 115.790 22.690 116.220 23.110 ;
        RECT 115.800 20.200 116.190 22.690 ;
        RECT 115.850 20.180 116.110 20.200 ;
      LAYER met3 ;
        RECT 16.800 220.470 17.120 220.510 ;
        RECT 26.000 220.470 26.460 221.220 ;
        RECT 16.800 220.170 26.460 220.470 ;
        RECT 16.800 220.130 17.120 220.170 ;
        RECT 26.000 220.100 26.460 220.170 ;
        RECT 77.620 213.735 78.430 217.675 ;
        RECT 42.665 209.110 45.155 209.135 ;
        RECT 77.710 209.120 78.370 213.735 ;
        RECT 114.990 209.120 117.360 209.165 ;
        RECT 47.110 209.110 117.360 209.120 ;
        RECT 9.070 206.535 12.260 209.085 ;
        RECT 19.220 206.855 25.350 208.815 ;
        RECT 42.660 206.620 117.360 209.110 ;
        RECT 42.660 206.610 45.740 206.620 ;
        RECT 42.665 206.585 45.155 206.610 ;
        RECT 114.990 205.645 117.360 206.620 ;
        RECT 125.090 182.525 128.090 182.570 ;
        RECT 125.070 181.385 129.510 182.525 ;
        RECT 0.950 174.490 8.390 174.950 ;
        RECT 125.090 174.490 128.090 181.385 ;
        RECT 0.950 171.490 128.180 174.490 ;
        RECT 0.950 170.590 8.390 171.490 ;
        RECT 0.960 30.385 5.130 33.865 ;
      LAYER met4 ;
        RECT 1.000 220.470 2.500 220.760 ;
        RECT 11.350 220.470 11.650 225.760 ;
        RECT 15.030 220.470 15.330 225.760 ;
        RECT 26.070 221.225 26.370 225.760 ;
        RECT 16.795 220.470 17.125 220.485 ;
        RECT 1.000 220.170 17.125 220.470 ;
        RECT 1.000 209.120 2.500 220.170 ;
        RECT 16.795 220.155 17.125 220.170 ;
        RECT 26.045 220.095 26.415 221.225 ;
        RECT 1.000 209.110 43.560 209.120 ;
        RECT 1.000 206.620 45.160 209.110 ;
        RECT 1.000 174.955 2.500 206.620 ;
        RECT 9.115 206.555 12.215 206.620 ;
        RECT 42.190 206.610 45.160 206.620 ;
        RECT 0.995 170.585 8.345 174.955 ;
        RECT 1.000 33.845 2.500 170.585 ;
        RECT 1.000 30.405 5.085 33.845 ;
        RECT 1.000 5.000 2.500 30.405 ;
    END
  END uio_oe[1]
  PIN uio_oe[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 7.670 224.760 7.970 225.760 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 3.990 224.760 4.290 225.760 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 59.190 224.760 59.490 225.760 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER li1 ;
        RECT 87.115 204.675 87.445 205.655 ;
        RECT 86.320 204.500 86.570 204.620 ;
        RECT 87.115 204.500 87.365 204.675 ;
        RECT 86.320 204.300 87.365 204.500 ;
        RECT 86.320 204.170 86.570 204.300 ;
        RECT 87.115 204.075 87.365 204.300 ;
        RECT 87.115 203.445 87.445 204.075 ;
      LAYER met1 ;
        RECT 84.560 204.710 85.280 206.210 ;
        RECT 85.430 204.900 86.370 204.930 ;
        RECT 85.430 204.710 86.590 204.900 ;
        RECT 84.560 204.680 86.590 204.710 ;
        RECT 84.560 204.110 86.600 204.680 ;
        RECT 84.560 203.930 86.590 204.110 ;
        RECT 84.560 203.730 85.430 203.930 ;
        RECT 85.590 203.900 86.590 203.930 ;
        RECT 84.590 203.710 85.430 203.730 ;
      LAYER met2 ;
        RECT 84.610 203.680 85.230 206.260 ;
      LAYER met3 ;
        RECT 60.970 222.530 61.290 222.550 ;
        RECT 60.920 222.510 61.290 222.530 ;
        RECT 64.300 222.510 64.680 222.520 ;
        RECT 60.920 222.210 64.680 222.510 ;
        RECT 60.920 222.170 61.290 222.210 ;
        RECT 64.300 222.200 64.680 222.210 ;
        RECT 60.920 222.150 61.240 222.170 ;
        RECT 84.560 203.705 85.280 206.235 ;
      LAYER met4 ;
        RECT 55.510 222.510 55.810 225.760 ;
        RECT 60.965 222.510 61.295 222.525 ;
        RECT 55.510 222.210 61.295 222.510 ;
        RECT 64.325 222.510 64.655 222.525 ;
        RECT 64.325 222.490 64.710 222.510 ;
        RECT 60.890 222.195 61.295 222.210 ;
        RECT 60.890 222.190 61.245 222.195 ;
        RECT 64.250 222.190 80.900 222.490 ;
        RECT 60.915 222.175 61.245 222.190 ;
        RECT 80.600 206.240 80.900 222.190 ;
        RECT 80.600 205.940 85.270 206.240 ;
        RECT 84.605 203.725 85.250 205.940 ;
        RECT 84.950 203.590 85.250 203.725 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 51.830 224.760 52.130 225.760 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 48.150 224.760 48.450 225.760 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER li1 ;
        RECT 58.325 219.475 58.655 220.255 ;
        RECT 57.890 219.455 58.655 219.475 ;
        RECT 59.165 219.455 59.495 220.255 ;
        RECT 57.890 219.285 59.495 219.455 ;
        RECT 57.890 219.280 58.155 219.285 ;
        RECT 57.650 218.800 58.155 219.280 ;
        RECT 57.890 218.695 58.155 218.800 ;
        RECT 57.890 218.515 59.495 218.695 ;
        RECT 58.325 218.045 58.655 218.515 ;
        RECT 59.165 218.045 59.495 218.515 ;
      LAYER met1 ;
        RECT 54.960 219.340 56.190 220.260 ;
        RECT 54.960 218.740 57.930 219.340 ;
        RECT 54.960 218.640 56.190 218.740 ;
        RECT 55.100 218.620 56.100 218.640 ;
      LAYER met2 ;
        RECT 55.010 218.590 56.140 220.310 ;
      LAYER met3 ;
        RECT 54.960 218.615 56.190 220.285 ;
      LAYER met4 ;
        RECT 44.470 221.670 44.770 225.760 ;
        RECT 44.390 221.370 55.840 221.670 ;
        RECT 55.540 220.265 55.840 221.370 ;
        RECT 55.005 218.635 56.145 220.265 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER li1 ;
        RECT 61.195 212.795 61.525 213.575 ;
        RECT 60.760 212.775 61.525 212.795 ;
        RECT 62.035 212.775 62.365 213.575 ;
        RECT 60.760 212.630 62.365 212.775 ;
        RECT 60.470 212.605 62.365 212.630 ;
        RECT 60.470 212.130 61.025 212.605 ;
        RECT 60.760 212.015 61.025 212.130 ;
        RECT 60.760 211.835 62.365 212.015 ;
        RECT 61.195 211.365 61.525 211.835 ;
        RECT 62.035 211.365 62.365 211.835 ;
      LAYER met1 ;
        RECT 54.160 212.870 55.660 212.890 ;
        RECT 54.160 212.690 56.100 212.870 ;
        RECT 54.160 212.090 56.150 212.690 ;
        RECT 59.440 212.090 60.820 212.690 ;
        RECT 54.160 211.870 56.100 212.090 ;
        RECT 60.010 212.070 60.820 212.090 ;
        RECT 54.160 211.840 55.660 211.870 ;
      LAYER met2 ;
        RECT 54.210 211.790 55.610 212.940 ;
        RECT 55.750 212.690 56.100 212.740 ;
        RECT 60.060 212.690 60.450 212.740 ;
        RECT 55.750 212.090 60.450 212.690 ;
        RECT 55.750 212.040 56.100 212.090 ;
        RECT 60.060 212.020 60.450 212.090 ;
      LAYER met3 ;
        RECT 54.160 211.815 55.660 212.915 ;
      LAYER met4 ;
        RECT 40.790 221.250 41.090 225.760 ;
        RECT 40.790 221.040 41.120 221.250 ;
        RECT 40.790 220.740 54.490 221.040 ;
        RECT 40.790 220.720 41.090 220.740 ;
        RECT 54.190 212.895 54.490 220.740 ;
        RECT 54.190 212.060 55.615 212.895 ;
        RECT 54.205 211.835 55.615 212.060 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 37.110 224.760 37.410 225.760 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 33.430 224.760 33.730 225.760 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.511500 ;
    PORT
      LAYER li1 ;
        RECT 98.575 194.005 98.910 195.435 ;
        RECT 98.855 190.730 99.170 191.155 ;
        RECT 98.855 190.715 99.320 190.730 ;
        RECT 98.855 190.465 99.545 190.715 ;
      LAYER met1 ;
        RECT 94.280 195.250 95.380 195.510 ;
        RECT 94.280 194.630 98.900 195.250 ;
        RECT 94.280 194.610 98.890 194.630 ;
        RECT 94.280 194.510 95.380 194.610 ;
        RECT 94.330 194.460 95.330 194.510 ;
        RECT 97.690 192.900 98.430 193.230 ;
        RECT 97.740 190.760 98.380 192.900 ;
        RECT 97.740 190.450 99.380 190.760 ;
      LAYER met2 ;
        RECT 94.330 194.460 95.330 195.560 ;
        RECT 97.750 193.280 98.380 195.010 ;
        RECT 97.740 192.850 98.380 193.280 ;
      LAYER met3 ;
        RECT 78.820 211.685 79.520 211.760 ;
        RECT 88.560 211.685 89.040 211.760 ;
        RECT 78.820 211.385 89.040 211.685 ;
        RECT 78.820 211.300 79.520 211.385 ;
        RECT 88.560 211.320 89.040 211.385 ;
        RECT 94.280 194.485 95.380 195.535 ;
      LAYER met4 ;
        RECT 88.630 211.760 88.930 225.760 ;
        RECT 78.875 211.350 79.205 211.680 ;
        RECT 78.890 195.360 79.190 211.350 ;
        RECT 88.560 211.320 89.040 211.760 ;
        RECT 94.325 195.360 95.335 195.515 ;
        RECT 78.890 195.060 95.335 195.360 ;
        RECT 94.180 194.870 95.335 195.060 ;
        RECT 94.325 194.505 95.335 194.870 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.511500 ;
    PORT
      LAYER li1 ;
        RECT 99.775 190.465 100.105 190.715 ;
        RECT 98.455 185.255 98.790 186.685 ;
      LAYER met1 ;
        RECT 99.750 190.140 100.120 190.720 ;
        RECT 99.690 189.870 100.170 190.140 ;
        RECT 93.370 186.620 94.620 186.630 ;
        RECT 93.370 186.490 94.630 186.620 ;
        RECT 93.370 186.460 94.840 186.490 ;
        RECT 98.470 186.470 98.780 186.480 ;
        RECT 93.370 185.830 95.130 186.460 ;
        RECT 97.040 185.840 98.780 186.470 ;
        RECT 98.470 185.830 98.780 185.840 ;
        RECT 93.370 185.800 94.840 185.830 ;
        RECT 93.370 185.630 94.630 185.800 ;
        RECT 93.630 185.620 94.630 185.630 ;
      LAYER met2 ;
        RECT 99.740 189.870 100.120 190.190 ;
        RECT 99.740 188.700 100.130 189.870 ;
        RECT 97.160 188.370 100.130 188.700 ;
        RECT 93.420 185.580 94.420 186.680 ;
        RECT 97.170 186.520 97.530 188.370 ;
        RECT 94.640 186.460 95.080 186.510 ;
        RECT 97.090 186.480 97.530 186.520 ;
        RECT 95.960 186.460 97.530 186.480 ;
        RECT 94.640 185.820 97.530 186.460 ;
        RECT 94.640 185.780 95.080 185.820 ;
        RECT 95.960 185.810 97.530 185.820 ;
        RECT 97.090 185.790 97.530 185.810 ;
      LAYER met3 ;
        RECT 79.740 210.960 80.180 211.050 ;
        RECT 84.860 210.960 85.300 210.980 ;
        RECT 79.740 210.660 85.300 210.960 ;
        RECT 79.740 210.570 80.180 210.660 ;
        RECT 84.860 210.500 85.300 210.660 ;
        RECT 79.700 193.680 80.270 196.770 ;
        RECT 79.730 193.670 80.250 193.680 ;
        RECT 93.370 185.605 94.620 186.655 ;
      LAYER met4 ;
        RECT 79.795 210.615 80.125 210.945 ;
        RECT 84.950 210.905 85.250 225.760 ;
        RECT 79.810 196.725 80.110 210.615 ;
        RECT 84.935 210.575 85.265 210.905 ;
        RECT 79.775 196.265 80.165 196.725 ;
        RECT 79.690 193.610 80.320 194.180 ;
        RECT 79.775 186.405 80.110 193.610 ;
        RECT 93.415 186.405 94.425 186.635 ;
        RECT 79.775 186.045 94.425 186.405 ;
        RECT 79.775 186.040 80.075 186.045 ;
        RECT 93.415 185.625 94.425 186.045 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER li1 ;
        RECT 134.495 203.550 135.330 203.620 ;
        RECT 134.495 203.540 135.765 203.550 ;
        RECT 133.650 203.430 135.765 203.540 ;
        RECT 133.650 203.385 134.625 203.430 ;
        RECT 133.650 203.210 134.575 203.385 ;
        RECT 135.205 203.375 135.765 203.430 ;
        RECT 135.245 203.220 135.765 203.375 ;
      LAYER met1 ;
        RECT 129.770 203.610 130.970 204.910 ;
        RECT 131.750 203.740 132.750 203.830 ;
        RECT 131.750 203.610 132.880 203.740 ;
        RECT 129.770 202.980 132.880 203.610 ;
        RECT 133.790 203.520 134.100 203.660 ;
        RECT 135.370 203.520 135.680 203.560 ;
        RECT 133.790 203.190 135.680 203.520 ;
        RECT 133.790 203.030 134.100 203.190 ;
        RECT 129.770 202.890 132.750 202.980 ;
        RECT 129.770 202.880 130.970 202.890 ;
        RECT 131.750 202.830 132.750 202.890 ;
      LAYER met2 ;
        RECT 129.820 202.830 130.920 204.960 ;
        RECT 132.420 203.580 132.930 203.690 ;
        RECT 133.740 203.580 134.150 203.610 ;
        RECT 132.420 203.110 134.150 203.580 ;
        RECT 132.420 203.030 132.930 203.110 ;
        RECT 133.740 203.080 134.150 203.110 ;
      LAYER met3 ;
        RECT 83.100 224.280 83.420 224.320 ;
        RECT 83.100 223.980 130.160 224.280 ;
        RECT 83.100 223.940 83.420 223.980 ;
        RECT 129.460 223.330 130.160 223.980 ;
        RECT 129.770 202.855 130.970 204.935 ;
      LAYER met4 ;
        RECT 81.270 224.280 81.570 225.760 ;
        RECT 83.095 224.280 83.425 224.295 ;
        RECT 81.270 223.980 83.425 224.280 ;
        RECT 83.095 223.965 83.425 223.980 ;
        RECT 129.505 223.325 130.115 224.285 ;
        RECT 129.810 204.915 130.110 223.325 ;
        RECT 129.810 204.100 130.925 204.915 ;
        RECT 129.815 202.875 130.925 204.100 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER li1 ;
        RECT 134.515 216.970 135.350 217.040 ;
        RECT 134.515 216.960 135.785 216.970 ;
        RECT 133.670 216.850 135.785 216.960 ;
        RECT 133.670 216.805 134.645 216.850 ;
        RECT 133.670 216.630 134.595 216.805 ;
        RECT 135.225 216.795 135.785 216.850 ;
        RECT 135.265 216.640 135.785 216.795 ;
      LAYER met1 ;
        RECT 128.380 217.060 129.300 217.130 ;
        RECT 131.750 217.120 132.750 217.220 ;
        RECT 131.750 217.060 132.920 217.120 ;
        RECT 128.380 216.360 132.920 217.060 ;
        RECT 133.830 216.980 134.140 217.070 ;
        RECT 133.830 216.610 135.690 216.980 ;
        RECT 133.830 216.600 135.450 216.610 ;
        RECT 133.830 216.440 134.140 216.600 ;
        RECT 128.380 216.300 132.750 216.360 ;
        RECT 128.380 216.230 129.300 216.300 ;
        RECT 131.750 216.220 132.750 216.300 ;
      LAYER met2 ;
        RECT 128.460 216.250 129.220 217.110 ;
        RECT 132.460 217.030 132.970 217.070 ;
        RECT 132.460 217.020 133.840 217.030 ;
        RECT 132.460 216.490 134.190 217.020 ;
        RECT 132.460 216.470 133.840 216.490 ;
        RECT 132.460 216.410 132.970 216.470 ;
      LAYER met3 ;
        RECT 79.370 223.450 79.690 223.490 ;
        RECT 128.140 223.450 128.810 223.460 ;
        RECT 79.370 223.150 128.810 223.450 ;
        RECT 79.370 223.110 79.690 223.150 ;
        RECT 128.140 222.390 128.810 223.150 ;
        RECT 128.410 216.275 129.270 217.085 ;
      LAYER met4 ;
        RECT 77.590 223.450 77.890 225.760 ;
        RECT 79.365 223.450 79.695 223.465 ;
        RECT 77.590 223.150 79.695 223.450 ;
        RECT 79.365 223.135 79.695 223.150 ;
        RECT 128.185 222.385 128.765 223.465 ;
        RECT 128.460 217.065 128.760 222.385 ;
        RECT 128.455 216.295 129.225 217.065 ;
        RECT 128.460 216.250 128.760 216.295 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER li1 ;
        RECT 30.120 213.210 30.450 213.645 ;
        RECT 30.120 213.125 30.520 213.210 ;
        RECT 30.275 213.085 30.520 213.125 ;
        RECT 30.330 212.505 30.520 213.085 ;
        RECT 30.285 212.455 30.520 212.505 ;
        RECT 30.110 212.375 30.520 212.455 ;
        RECT 30.110 211.530 30.440 212.375 ;
      LAYER met1 ;
        RECT 45.430 223.360 48.390 223.680 ;
        RECT 45.480 216.490 45.780 223.360 ;
        RECT 44.340 215.950 45.840 216.490 ;
        RECT 30.900 214.720 31.670 215.430 ;
        RECT 30.030 214.340 31.670 214.720 ;
        RECT 30.540 214.330 31.670 214.340 ;
        RECT 30.090 213.550 30.420 213.560 ;
        RECT 30.060 213.170 30.510 213.550 ;
      LAYER met2 ;
        RECT 45.480 223.310 48.340 223.730 ;
        RECT 44.390 215.900 45.790 216.540 ;
        RECT 30.080 214.290 30.510 214.770 ;
        RECT 30.110 213.570 30.470 214.290 ;
        RECT 30.950 214.280 31.620 215.480 ;
        RECT 30.110 213.120 30.460 213.570 ;
      LAYER met3 ;
        RECT 71.610 223.760 74.290 223.920 ;
        RECT 45.380 223.460 74.290 223.760 ;
        RECT 45.430 223.335 48.390 223.460 ;
        RECT 44.340 216.250 45.840 216.515 ;
        RECT 31.130 215.950 45.840 216.250 ;
        RECT 31.130 215.455 31.430 215.950 ;
        RECT 44.340 215.925 45.840 215.950 ;
        RECT 30.900 214.305 31.670 215.455 ;
      LAYER met4 ;
        RECT 73.910 223.870 74.210 225.760 ;
        RECT 71.690 223.410 74.260 223.870 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER li1 ;
        RECT 42.030 213.210 42.360 213.645 ;
        RECT 42.030 213.125 42.430 213.210 ;
        RECT 42.185 213.085 42.430 213.125 ;
        RECT 42.240 212.505 42.430 213.085 ;
        RECT 42.195 212.455 42.430 212.505 ;
        RECT 42.020 212.375 42.430 212.455 ;
        RECT 42.020 211.530 42.350 212.375 ;
      LAYER met1 ;
        RECT 42.070 223.290 43.670 224.310 ;
        RECT 41.910 214.800 42.970 214.810 ;
        RECT 43.110 214.800 43.410 223.290 ;
        RECT 41.910 214.460 43.410 214.800 ;
        RECT 42.850 214.390 43.410 214.460 ;
        RECT 42.850 214.380 43.400 214.390 ;
        RECT 41.990 213.560 42.320 213.570 ;
        RECT 41.970 213.230 42.410 213.560 ;
      LAYER met2 ;
        RECT 42.120 223.240 43.620 224.360 ;
        RECT 41.960 214.410 42.430 214.860 ;
        RECT 42.010 213.580 42.360 214.410 ;
        RECT 42.020 213.180 42.360 213.580 ;
      LAYER met3 ;
        RECT 68.180 224.370 70.570 224.620 ;
        RECT 42.060 224.120 70.570 224.370 ;
        RECT 42.060 224.070 70.550 224.120 ;
        RECT 42.070 223.265 43.670 224.070 ;
      LAYER met4 ;
        RECT 70.230 224.625 70.530 225.760 ;
        RECT 68.225 224.440 70.530 224.625 ;
        RECT 68.225 224.115 70.525 224.440 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER li1 ;
        RECT 30.450 201.235 30.780 202.080 ;
        RECT 30.450 201.155 30.860 201.235 ;
        RECT 30.625 201.105 30.860 201.155 ;
        RECT 30.670 200.525 30.860 201.105 ;
        RECT 30.615 200.485 30.860 200.525 ;
        RECT 30.460 200.400 30.860 200.485 ;
        RECT 30.460 199.965 30.790 200.400 ;
      LAYER met1 ;
        RECT 46.860 214.750 47.430 217.620 ;
        RECT 46.960 205.790 47.260 214.750 ;
        RECT 30.960 205.490 47.260 205.790 ;
        RECT 30.960 203.790 31.260 205.490 ;
        RECT 30.560 202.790 31.560 203.790 ;
        RECT 30.410 200.080 31.280 200.350 ;
      LAYER met2 ;
        RECT 46.520 222.570 50.740 223.020 ;
        RECT 46.970 217.670 47.270 222.570 ;
        RECT 46.910 214.700 47.380 217.670 ;
        RECT 30.830 203.380 31.170 203.410 ;
        RECT 30.810 200.400 31.170 203.380 ;
        RECT 30.810 200.030 31.230 200.400 ;
      LAYER met3 ;
        RECT 50.740 223.060 67.420 223.160 ;
        RECT 50.460 222.995 67.420 223.060 ;
        RECT 46.470 222.860 67.420 222.995 ;
        RECT 46.470 222.595 51.450 222.860 ;
        RECT 65.130 222.840 67.420 222.860 ;
        RECT 50.460 222.560 51.450 222.595 ;
      LAYER met4 ;
        RECT 66.550 223.165 66.850 225.760 ;
        RECT 65.175 222.835 67.375 223.165 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER li1 ;
        RECT 42.770 201.215 43.100 202.060 ;
        RECT 42.770 201.135 43.180 201.215 ;
        RECT 42.945 201.085 43.180 201.135 ;
        RECT 42.990 200.505 43.180 201.085 ;
        RECT 42.935 200.465 43.180 200.505 ;
        RECT 42.780 200.380 43.180 200.465 ;
        RECT 42.780 199.945 43.110 200.380 ;
      LAYER met1 ;
        RECT 51.920 221.060 63.400 221.360 ;
        RECT 52.220 203.830 52.760 221.060 ;
        RECT 60.740 221.040 63.400 221.060 ;
        RECT 60.750 220.890 63.300 221.040 ;
        RECT 42.940 203.290 52.760 203.830 ;
        RECT 42.940 202.830 43.940 203.290 ;
        RECT 42.720 200.060 43.660 200.360 ;
      LAYER met2 ;
        RECT 60.840 220.840 63.250 221.260 ;
        RECT 43.090 202.810 43.720 203.340 ;
        RECT 43.150 200.070 43.720 202.810 ;
        RECT 43.160 200.010 43.610 200.070 ;
      LAYER met3 ;
        RECT 60.790 220.865 63.300 221.235 ;
      LAYER met4 ;
        RECT 62.870 221.215 63.170 225.760 ;
        RECT 60.835 220.885 63.255 221.215 ;
        RECT 62.870 220.830 63.170 220.885 ;
    END
  END uo_out[7]
  OBS
      LAYER pwell ;
        RECT 57.815 217.895 60.005 218.805 ;
        RECT 60.495 217.895 62.685 218.805 ;
        RECT 63.175 217.895 65.365 218.805 ;
        RECT 65.910 218.575 68.190 218.805 ;
        RECT 71.395 218.575 72.325 218.795 ;
        RECT 65.910 217.895 76.835 218.575 ;
        RECT 59.745 217.705 59.915 217.895 ;
        RECT 62.425 217.705 62.595 217.895 ;
        RECT 65.105 217.705 65.275 217.895 ;
        RECT 76.525 217.705 76.695 217.895 ;
        RECT 66.775 214.555 68.965 215.465 ;
        RECT 66.865 214.365 67.035 214.555 ;
        RECT 10.565 213.835 10.735 214.025 ;
        RECT 23.365 213.845 23.535 214.035 ;
        RECT 35.275 213.845 35.445 214.035 ;
        RECT 10.425 213.155 19.155 213.835 ;
        RECT 23.225 213.165 31.955 213.845 ;
        RECT 35.135 213.165 43.865 213.845 ;
        RECT 13.940 212.935 14.850 213.155 ;
        RECT 16.390 212.925 19.155 213.155 ;
        RECT 26.740 212.945 27.650 213.165 ;
        RECT 29.190 212.935 31.955 213.165 ;
        RECT 38.650 212.945 39.560 213.165 ;
        RECT 41.100 212.935 43.865 213.165 ;
        RECT 60.685 211.215 62.875 212.125 ;
        RECT 63.365 211.215 65.555 212.125 ;
        RECT 65.910 211.895 68.190 212.125 ;
        RECT 71.395 211.895 72.325 212.115 ;
        RECT 65.910 211.215 76.835 211.895 ;
        RECT 62.615 211.025 62.785 211.215 ;
        RECT 65.295 211.025 65.465 211.215 ;
        RECT 76.525 211.025 76.695 211.215 ;
        RECT 86.605 203.295 87.955 204.205 ;
        RECT 88.175 203.295 89.525 204.205 ;
        RECT 89.775 203.975 92.540 204.205 ;
        RECT 94.080 203.975 94.990 204.195 ;
        RECT 98.685 203.975 101.450 204.205 ;
        RECT 102.990 203.975 103.900 204.195 ;
        RECT 107.595 203.975 110.360 204.205 ;
        RECT 111.900 203.975 112.810 204.195 ;
        RECT 89.775 203.295 98.505 203.975 ;
        RECT 98.685 203.295 107.415 203.975 ;
        RECT 107.595 203.295 116.325 203.975 ;
        RECT 87.655 203.105 87.825 203.295 ;
        RECT 89.225 203.105 89.395 203.295 ;
        RECT 98.195 203.105 98.365 203.295 ;
        RECT 107.105 203.105 107.275 203.295 ;
        RECT 116.015 203.105 116.185 203.295 ;
        RECT 103.445 189.475 105.635 190.385 ;
        RECT 103.535 189.285 103.705 189.475 ;
      LAYER li1 ;
        RECT 61.005 219.475 61.335 220.255 ;
        RECT 60.570 219.455 61.335 219.475 ;
        RECT 61.845 219.455 62.175 220.255 ;
        RECT 63.685 219.475 64.015 220.255 ;
        RECT 60.570 219.285 62.175 219.455 ;
        RECT 63.250 219.455 64.015 219.475 ;
        RECT 64.525 219.455 64.855 220.255 ;
        RECT 63.250 219.285 64.855 219.455 ;
        RECT 66.420 219.870 66.720 220.255 ;
        RECT 66.420 219.325 66.810 219.870 ;
        RECT 68.280 219.825 68.505 220.255 ;
        RECT 69.310 219.875 69.480 220.165 ;
        RECT 67.005 219.655 68.505 219.825 ;
        RECT 58.325 219.110 59.955 219.115 ;
        RECT 60.570 219.110 60.835 219.285 ;
        RECT 58.325 218.880 60.835 219.110 ;
        RECT 58.325 218.865 59.955 218.880 ;
        RECT 60.570 218.695 60.835 218.880 ;
        RECT 61.005 219.110 62.635 219.115 ;
        RECT 63.250 219.110 63.515 219.285 ;
        RECT 61.005 218.880 63.515 219.110 ;
        RECT 61.005 218.865 62.635 218.880 ;
        RECT 63.250 218.695 63.515 218.880 ;
        RECT 63.685 218.865 65.315 219.115 ;
        RECT 60.570 218.515 62.175 218.695 ;
        RECT 63.250 218.515 64.855 218.695 ;
        RECT 61.005 218.045 61.335 218.515 ;
        RECT 61.845 218.045 62.175 218.515 ;
        RECT 63.685 218.045 64.015 218.515 ;
        RECT 64.525 218.045 64.855 218.515 ;
        RECT 66.420 218.615 66.590 219.325 ;
        RECT 67.005 219.115 67.175 219.655 ;
        RECT 67.850 219.585 68.505 219.655 ;
        RECT 68.680 219.705 69.480 219.875 ;
        RECT 70.070 219.915 70.940 220.255 ;
        RECT 66.760 218.785 67.175 219.115 ;
        RECT 66.420 218.100 66.800 218.615 ;
        RECT 67.345 218.055 67.680 219.485 ;
        RECT 67.850 218.675 68.020 219.585 ;
        RECT 68.680 219.115 68.850 219.705 ;
        RECT 70.070 219.535 70.240 219.915 ;
        RECT 71.175 219.795 71.345 220.255 ;
        RECT 72.180 219.825 72.350 220.165 ;
        RECT 73.085 219.825 73.255 220.165 ;
        RECT 69.020 219.365 70.240 219.535 ;
        RECT 70.410 219.455 70.870 219.745 ;
        RECT 71.175 219.625 71.735 219.795 ;
        RECT 72.180 219.655 73.255 219.825 ;
        RECT 73.425 219.925 74.105 220.255 ;
        RECT 74.320 219.925 74.570 220.255 ;
        RECT 71.565 219.485 71.735 219.625 ;
        RECT 70.410 219.445 71.375 219.455 ;
        RECT 70.070 219.275 70.240 219.365 ;
        RECT 70.700 219.285 71.375 219.445 ;
        RECT 68.190 219.085 68.850 219.115 ;
        RECT 68.190 218.865 69.025 219.085 ;
        RECT 68.680 218.785 69.025 218.865 ;
        RECT 67.850 218.505 68.505 218.675 ;
        RECT 68.255 218.135 68.505 218.505 ;
        RECT 68.855 218.255 69.025 218.785 ;
        RECT 69.195 218.825 69.735 219.195 ;
        RECT 70.070 219.105 70.475 219.275 ;
        RECT 69.195 218.425 69.435 218.825 ;
        RECT 69.915 218.655 70.135 218.935 ;
        RECT 69.605 218.485 70.135 218.655 ;
        RECT 69.605 218.255 69.775 218.485 ;
        RECT 68.855 218.085 69.775 218.255 ;
        RECT 70.305 218.325 70.475 219.105 ;
        RECT 70.645 218.495 70.995 219.115 ;
        RECT 71.165 218.495 71.375 219.285 ;
        RECT 71.565 219.315 73.065 219.485 ;
        RECT 71.565 218.625 71.735 219.315 ;
        RECT 73.425 219.145 73.595 219.925 ;
        RECT 74.400 219.795 74.570 219.925 ;
        RECT 71.905 218.975 73.595 219.145 ;
        RECT 73.765 219.365 74.230 219.755 ;
        RECT 74.400 219.625 74.795 219.795 ;
        RECT 71.905 218.795 72.075 218.975 ;
        RECT 70.305 218.045 71.255 218.325 ;
        RECT 71.565 218.235 71.825 218.625 ;
        RECT 72.245 218.555 73.035 218.805 ;
        RECT 71.475 218.065 71.825 218.235 ;
        RECT 73.240 218.265 73.410 218.975 ;
        RECT 73.765 218.775 73.935 219.365 ;
        RECT 73.580 218.555 73.935 218.775 ;
        RECT 74.105 218.555 74.455 219.175 ;
        RECT 74.625 218.265 74.795 219.625 ;
        RECT 73.240 218.095 74.095 218.265 ;
        RECT 74.300 218.095 74.795 218.265 ;
        RECT 75.655 218.135 75.825 220.255 ;
        RECT 76.495 219.755 76.750 220.255 ;
        RECT 76.000 219.585 76.750 219.755 ;
        RECT 76.000 218.595 76.230 219.585 ;
        RECT 133.625 218.670 135.825 218.885 ;
        RECT 76.000 218.425 76.750 218.595 ;
        RECT 133.625 218.550 134.595 218.670 ;
        RECT 135.205 218.630 135.825 218.670 ;
        RECT 76.495 218.135 76.750 218.425 ;
        RECT 134.765 217.975 135.095 218.500 ;
        RECT 133.645 217.905 135.095 217.975 ;
        RECT 133.645 217.705 135.745 217.905 ;
        RECT 133.645 217.645 134.375 217.705 ;
        RECT 135.475 217.645 135.745 217.705 ;
        RECT 63.665 215.775 63.980 216.215 ;
        RECT 64.315 216.195 64.615 216.745 ;
        RECT 65.345 216.365 65.795 216.915 ;
        RECT 64.315 216.025 65.255 216.195 ;
        RECT 65.085 215.775 65.255 216.025 ;
        RECT 63.665 215.525 64.355 215.775 ;
        RECT 64.585 215.525 64.915 215.775 ;
        RECT 65.085 215.445 65.375 215.775 ;
        RECT 65.545 215.770 65.795 216.365 ;
        RECT 67.285 216.115 67.615 216.915 ;
        RECT 68.125 216.135 68.455 216.915 ;
        RECT 68.125 216.115 68.890 216.135 ;
        RECT 134.765 216.130 135.095 216.680 ;
        RECT 134.765 216.120 135.790 216.130 ;
        RECT 67.285 215.945 68.890 216.115 ;
        RECT 66.825 215.770 68.455 215.775 ;
        RECT 65.545 215.525 68.455 215.770 ;
        RECT 65.545 215.520 66.830 215.525 ;
        RECT 65.085 215.355 65.255 215.445 ;
        RECT 63.865 215.165 65.255 215.355 ;
        RECT 63.865 214.805 64.195 215.165 ;
        RECT 65.545 214.995 65.795 215.520 ;
        RECT 68.625 215.355 68.890 215.945 ;
        RECT 133.625 215.930 135.790 216.120 ;
        RECT 133.625 215.780 134.560 215.930 ;
        RECT 135.265 215.800 135.790 215.930 ;
        RECT 65.245 214.705 65.795 214.995 ;
        RECT 67.285 215.175 68.890 215.355 ;
        RECT 134.185 215.220 134.560 215.780 ;
        RECT 67.285 214.705 67.615 215.175 ;
        RECT 68.125 214.705 68.455 215.175 ;
        RECT 134.765 215.050 135.095 215.760 ;
        RECT 133.755 214.880 135.725 215.050 ;
        RECT 133.755 214.165 133.925 214.880 ;
        RECT 134.095 214.390 135.385 214.710 ;
        RECT 135.055 214.245 135.385 214.390 ;
        RECT 135.555 214.265 135.725 214.880 ;
        RECT 134.125 214.030 134.845 214.220 ;
        RECT 133.625 213.860 133.955 213.940 ;
        RECT 135.555 213.860 135.725 214.095 ;
        RECT 10.595 213.305 10.765 213.595 ;
        RECT 10.595 213.135 11.260 213.305 ;
        RECT 11.030 212.145 11.260 213.135 ;
        RECT 10.595 211.975 11.260 212.145 ;
        RECT 10.595 211.475 10.765 211.975 ;
        RECT 11.435 211.475 11.620 213.595 ;
        RECT 12.295 213.405 12.630 213.575 ;
        RECT 12.825 213.405 13.500 213.575 ;
        RECT 12.295 213.265 12.465 213.405 ;
        RECT 11.790 212.275 12.070 213.225 ;
        RECT 12.240 213.135 12.465 213.265 ;
        RECT 12.240 212.030 12.410 213.135 ;
        RECT 12.635 212.985 13.160 213.205 ;
        RECT 12.580 212.220 12.820 212.815 ;
        RECT 12.990 212.285 13.160 212.985 ;
        RECT 13.330 212.625 13.500 213.405 ;
        RECT 14.370 213.405 14.775 213.575 ;
        RECT 14.945 213.405 15.730 213.575 ;
        RECT 14.370 213.175 14.540 213.405 ;
        RECT 13.710 212.875 14.540 213.175 ;
        RECT 14.925 212.905 15.390 213.235 ;
        RECT 13.710 212.845 13.910 212.875 ;
        RECT 14.030 212.625 14.200 212.695 ;
        RECT 13.330 212.455 14.200 212.625 ;
        RECT 13.690 212.365 14.200 212.455 ;
        RECT 12.240 211.900 12.545 212.030 ;
        RECT 12.990 211.920 13.520 212.285 ;
        RECT 12.295 211.475 12.545 211.900 ;
        RECT 13.690 211.750 13.860 212.365 ;
        RECT 12.755 211.580 13.860 211.750 ;
        RECT 14.370 211.805 14.540 212.875 ;
        RECT 14.710 211.975 14.900 212.695 ;
        RECT 15.070 211.945 15.390 212.905 ;
        RECT 15.560 212.945 15.730 213.405 ;
        RECT 16.480 213.115 16.810 213.640 ;
        RECT 17.320 213.200 17.650 213.635 ;
        RECT 17.840 213.325 18.090 213.595 ;
        RECT 17.320 213.115 17.720 213.200 ;
        RECT 16.610 212.945 16.810 213.115 ;
        RECT 17.475 213.075 17.720 213.115 ;
        RECT 15.560 212.615 16.440 212.945 ;
        RECT 16.610 212.615 17.360 212.945 ;
        RECT 14.370 211.475 14.620 211.805 ;
        RECT 15.560 211.775 15.730 212.615 ;
        RECT 16.610 212.410 16.800 212.615 ;
        RECT 17.530 212.495 17.720 213.075 ;
        RECT 17.485 212.445 17.720 212.495 ;
        RECT 15.900 212.035 16.800 212.410 ;
        RECT 14.845 211.605 15.730 211.775 ;
        RECT 16.460 211.475 16.800 212.035 ;
        RECT 17.310 212.365 17.720 212.445 ;
        RECT 17.890 212.945 18.090 213.325 ;
        RECT 18.815 213.030 19.070 213.685 ;
        RECT 23.395 213.315 23.565 213.605 ;
        RECT 23.395 213.145 24.060 213.315 ;
        RECT 17.890 212.615 18.665 212.945 ;
        RECT 17.310 211.520 17.640 212.365 ;
        RECT 17.890 212.225 18.160 212.615 ;
        RECT 18.835 212.460 19.070 213.030 ;
        RECT 17.830 211.495 18.160 212.225 ;
        RECT 18.735 211.475 19.070 212.460 ;
        RECT 23.310 212.325 23.660 212.975 ;
        RECT 23.830 212.155 24.060 213.145 ;
        RECT 23.395 211.985 24.060 212.155 ;
        RECT 23.395 211.485 23.565 211.985 ;
        RECT 24.235 211.485 24.420 213.605 ;
        RECT 25.095 213.415 25.430 213.585 ;
        RECT 25.625 213.415 26.300 213.585 ;
        RECT 25.095 213.275 25.265 213.415 ;
        RECT 24.590 212.285 24.870 213.235 ;
        RECT 25.040 213.145 25.265 213.275 ;
        RECT 25.040 212.040 25.210 213.145 ;
        RECT 25.435 212.995 25.960 213.215 ;
        RECT 25.380 212.230 25.620 212.825 ;
        RECT 25.790 212.295 25.960 212.995 ;
        RECT 26.130 212.635 26.300 213.415 ;
        RECT 27.170 213.415 27.575 213.585 ;
        RECT 27.745 213.415 28.530 213.585 ;
        RECT 27.170 213.185 27.340 213.415 ;
        RECT 26.510 212.885 27.340 213.185 ;
        RECT 27.725 212.915 28.190 213.245 ;
        RECT 26.510 212.855 26.710 212.885 ;
        RECT 26.830 212.635 27.000 212.705 ;
        RECT 26.130 212.465 27.000 212.635 ;
        RECT 26.490 212.375 27.000 212.465 ;
        RECT 25.040 211.910 25.345 212.040 ;
        RECT 25.790 211.930 26.320 212.295 ;
        RECT 25.095 211.485 25.345 211.910 ;
        RECT 26.490 211.760 26.660 212.375 ;
        RECT 25.555 211.590 26.660 211.760 ;
        RECT 27.170 211.815 27.340 212.885 ;
        RECT 27.510 211.985 27.700 212.705 ;
        RECT 27.870 211.955 28.190 212.915 ;
        RECT 28.360 212.955 28.530 213.415 ;
        RECT 29.280 213.125 29.610 213.650 ;
        RECT 30.640 213.335 30.890 213.605 ;
        RECT 29.410 212.955 29.610 213.125 ;
        RECT 30.690 212.955 30.890 213.335 ;
        RECT 31.615 213.040 31.870 213.695 ;
        RECT 35.305 213.315 35.475 213.605 ;
        RECT 35.305 213.145 35.970 213.315 ;
        RECT 28.360 212.625 29.240 212.955 ;
        RECT 29.410 212.625 30.160 212.955 ;
        RECT 30.690 212.625 31.465 212.955 ;
        RECT 27.170 211.485 27.420 211.815 ;
        RECT 28.360 211.785 28.530 212.625 ;
        RECT 29.410 212.420 29.600 212.625 ;
        RECT 28.700 212.045 29.600 212.420 ;
        RECT 30.690 212.235 30.960 212.625 ;
        RECT 31.635 212.470 31.870 213.040 ;
        RECT 35.220 212.890 35.570 212.975 ;
        RECT 35.210 212.630 35.570 212.890 ;
        RECT 27.645 211.615 28.530 211.785 ;
        RECT 29.260 211.485 29.600 212.045 ;
        RECT 30.630 211.505 30.960 212.235 ;
        RECT 31.535 211.485 31.870 212.470 ;
        RECT 35.220 212.325 35.570 212.630 ;
        RECT 35.740 212.155 35.970 213.145 ;
        RECT 35.305 211.985 35.970 212.155 ;
        RECT 35.305 211.485 35.475 211.985 ;
        RECT 36.145 211.485 36.330 213.605 ;
        RECT 37.005 213.415 37.340 213.585 ;
        RECT 37.535 213.415 38.210 213.585 ;
        RECT 37.005 213.275 37.175 213.415 ;
        RECT 36.500 212.285 36.780 213.235 ;
        RECT 36.950 213.145 37.175 213.275 ;
        RECT 36.950 212.040 37.120 213.145 ;
        RECT 37.345 212.995 37.870 213.215 ;
        RECT 37.290 212.230 37.530 212.825 ;
        RECT 37.700 212.295 37.870 212.995 ;
        RECT 38.040 212.635 38.210 213.415 ;
        RECT 39.080 213.415 39.485 213.585 ;
        RECT 39.655 213.415 40.440 213.585 ;
        RECT 39.080 213.185 39.250 213.415 ;
        RECT 38.420 212.885 39.250 213.185 ;
        RECT 39.635 212.915 40.100 213.245 ;
        RECT 38.420 212.855 38.620 212.885 ;
        RECT 38.740 212.635 38.910 212.705 ;
        RECT 38.040 212.465 38.910 212.635 ;
        RECT 38.400 212.375 38.910 212.465 ;
        RECT 36.950 211.910 37.255 212.040 ;
        RECT 37.700 211.930 38.230 212.295 ;
        RECT 37.005 211.485 37.255 211.910 ;
        RECT 38.400 211.760 38.570 212.375 ;
        RECT 37.465 211.590 38.570 211.760 ;
        RECT 39.080 211.815 39.250 212.885 ;
        RECT 39.420 211.985 39.610 212.705 ;
        RECT 39.780 211.955 40.100 212.915 ;
        RECT 40.270 212.955 40.440 213.415 ;
        RECT 41.190 213.125 41.520 213.650 ;
        RECT 42.550 213.335 42.800 213.605 ;
        RECT 41.320 212.955 41.520 213.125 ;
        RECT 42.600 212.955 42.800 213.335 ;
        RECT 43.525 213.040 43.780 213.695 ;
        RECT 133.625 213.690 135.725 213.860 ;
        RECT 40.270 212.625 41.150 212.955 ;
        RECT 41.320 212.625 42.070 212.955 ;
        RECT 42.600 212.625 43.375 212.955 ;
        RECT 39.080 211.485 39.330 211.815 ;
        RECT 40.270 211.785 40.440 212.625 ;
        RECT 41.320 212.420 41.510 212.625 ;
        RECT 40.610 212.045 41.510 212.420 ;
        RECT 42.600 212.235 42.870 212.625 ;
        RECT 43.545 212.470 43.780 213.040 ;
        RECT 63.875 212.795 64.205 213.575 ;
        RECT 39.555 211.615 40.440 211.785 ;
        RECT 41.170 211.485 41.510 212.045 ;
        RECT 42.540 211.505 42.870 212.235 ;
        RECT 43.445 211.485 43.780 212.470 ;
        RECT 63.440 212.775 64.205 212.795 ;
        RECT 64.715 212.775 65.045 213.575 ;
        RECT 63.440 212.605 65.045 212.775 ;
        RECT 66.420 213.190 66.720 213.575 ;
        RECT 66.420 212.645 66.810 213.190 ;
        RECT 68.280 213.145 68.505 213.575 ;
        RECT 69.310 213.195 69.480 213.485 ;
        RECT 67.005 212.975 68.505 213.145 ;
        RECT 61.195 212.430 62.825 212.435 ;
        RECT 63.440 212.430 63.705 212.605 ;
        RECT 61.195 212.190 63.705 212.430 ;
        RECT 61.195 212.185 62.825 212.190 ;
        RECT 63.440 212.015 63.705 212.190 ;
        RECT 63.875 212.185 65.505 212.435 ;
        RECT 63.440 211.835 65.045 212.015 ;
        RECT 63.875 211.365 64.205 211.835 ;
        RECT 64.715 211.365 65.045 211.835 ;
        RECT 66.420 211.935 66.590 212.645 ;
        RECT 67.005 212.435 67.175 212.975 ;
        RECT 67.850 212.905 68.505 212.975 ;
        RECT 68.680 213.025 69.480 213.195 ;
        RECT 70.070 213.235 70.940 213.575 ;
        RECT 66.760 212.105 67.175 212.435 ;
        RECT 66.420 211.420 66.800 211.935 ;
        RECT 67.345 211.375 67.680 212.805 ;
        RECT 67.850 211.995 68.020 212.905 ;
        RECT 68.680 212.435 68.850 213.025 ;
        RECT 70.070 212.855 70.240 213.235 ;
        RECT 71.175 213.115 71.345 213.575 ;
        RECT 72.180 213.145 72.350 213.485 ;
        RECT 73.085 213.145 73.255 213.485 ;
        RECT 69.020 212.685 70.240 212.855 ;
        RECT 70.410 212.775 70.870 213.065 ;
        RECT 71.175 212.945 71.735 213.115 ;
        RECT 72.180 212.975 73.255 213.145 ;
        RECT 73.425 213.245 74.105 213.575 ;
        RECT 74.320 213.245 74.570 213.575 ;
        RECT 71.565 212.805 71.735 212.945 ;
        RECT 70.410 212.765 71.375 212.775 ;
        RECT 70.070 212.595 70.240 212.685 ;
        RECT 70.700 212.605 71.375 212.765 ;
        RECT 68.190 212.405 68.850 212.435 ;
        RECT 68.190 212.185 69.025 212.405 ;
        RECT 68.680 212.105 69.025 212.185 ;
        RECT 67.850 211.825 68.505 211.995 ;
        RECT 68.255 211.455 68.505 211.825 ;
        RECT 68.855 211.575 69.025 212.105 ;
        RECT 69.195 212.145 69.735 212.515 ;
        RECT 70.070 212.425 70.475 212.595 ;
        RECT 69.195 211.745 69.435 212.145 ;
        RECT 69.915 211.975 70.135 212.255 ;
        RECT 69.605 211.805 70.135 211.975 ;
        RECT 69.605 211.575 69.775 211.805 ;
        RECT 68.855 211.405 69.775 211.575 ;
        RECT 70.305 211.645 70.475 212.425 ;
        RECT 70.645 211.815 70.995 212.435 ;
        RECT 71.165 211.815 71.375 212.605 ;
        RECT 71.565 212.635 73.065 212.805 ;
        RECT 71.565 211.945 71.735 212.635 ;
        RECT 73.425 212.465 73.595 213.245 ;
        RECT 74.400 213.115 74.570 213.245 ;
        RECT 71.905 212.295 73.595 212.465 ;
        RECT 73.765 212.685 74.230 213.075 ;
        RECT 74.400 212.945 74.795 213.115 ;
        RECT 71.905 212.115 72.075 212.295 ;
        RECT 70.305 211.365 71.255 211.645 ;
        RECT 71.565 211.555 71.825 211.945 ;
        RECT 72.245 211.875 73.035 212.125 ;
        RECT 71.475 211.385 71.825 211.555 ;
        RECT 73.240 211.585 73.410 212.295 ;
        RECT 73.765 212.095 73.935 212.685 ;
        RECT 73.580 211.875 73.935 212.095 ;
        RECT 74.105 211.875 74.455 212.495 ;
        RECT 74.625 211.585 74.795 212.945 ;
        RECT 73.240 211.415 74.095 211.585 ;
        RECT 74.300 211.415 74.795 211.585 ;
        RECT 75.655 211.455 75.825 213.575 ;
        RECT 76.495 213.075 76.750 213.575 ;
        RECT 134.515 213.350 134.845 213.520 ;
        RECT 134.515 213.180 134.775 213.350 ;
        RECT 135.025 213.230 135.325 213.690 ;
        RECT 76.000 212.905 76.750 213.075 ;
        RECT 133.730 213.010 134.775 213.180 ;
        RECT 134.995 213.030 135.325 213.230 ;
        RECT 76.000 211.915 76.230 212.905 ;
        RECT 133.730 212.075 133.900 213.010 ;
        RECT 134.070 212.480 134.435 212.840 ;
        RECT 134.605 212.820 134.775 213.010 ;
        RECT 134.605 212.650 135.725 212.820 ;
        RECT 134.070 212.310 135.355 212.480 ;
        RECT 76.000 211.745 76.750 211.915 ;
        RECT 134.370 211.900 134.965 212.140 ;
        RECT 135.135 211.955 135.355 212.310 ;
        RECT 135.555 212.145 135.725 212.650 ;
        RECT 76.495 211.455 76.750 211.745 ;
        RECT 133.625 211.730 134.180 211.865 ;
        RECT 135.555 211.785 135.725 211.950 ;
        RECT 135.285 211.730 135.725 211.785 ;
        RECT 133.625 211.615 135.725 211.730 ;
        RECT 134.050 211.560 135.415 211.615 ;
        RECT 134.425 211.110 135.375 211.390 ;
        RECT 133.625 210.755 135.745 210.940 ;
        RECT 134.125 210.350 135.455 210.580 ;
        RECT 134.125 210.085 134.295 210.350 ;
        RECT 133.625 209.915 134.295 210.085 ;
        RECT 134.465 209.830 135.115 210.180 ;
        RECT 135.285 210.085 135.455 210.350 ;
        RECT 135.285 209.915 135.745 210.085 ;
        RECT 88.685 204.675 89.015 205.655 ;
        RECT 87.535 204.510 87.865 204.515 ;
        RECT 88.685 204.510 88.935 204.675 ;
        RECT 89.860 204.670 90.195 205.655 ;
        RECT 90.770 204.905 91.100 205.635 ;
        RECT 87.535 204.270 88.935 204.510 ;
        RECT 87.535 204.265 87.865 204.270 ;
        RECT 88.685 204.075 88.935 204.270 ;
        RECT 89.105 204.265 89.435 204.515 ;
        RECT 89.860 204.100 90.095 204.670 ;
        RECT 90.770 204.515 91.040 204.905 ;
        RECT 91.290 204.765 91.620 205.610 ;
        RECT 90.265 204.185 91.040 204.515 ;
        RECT 88.685 203.445 89.015 204.075 ;
        RECT 89.860 203.445 90.115 204.100 ;
        RECT 90.840 203.805 91.040 204.185 ;
        RECT 91.210 204.685 91.620 204.765 ;
        RECT 92.130 205.095 92.470 205.655 ;
        RECT 93.200 205.355 94.085 205.525 ;
        RECT 92.130 204.720 93.030 205.095 ;
        RECT 91.210 204.635 91.445 204.685 ;
        RECT 91.210 204.055 91.400 204.635 ;
        RECT 92.130 204.515 92.320 204.720 ;
        RECT 93.200 204.515 93.370 205.355 ;
        RECT 94.310 205.325 94.560 205.655 ;
        RECT 91.570 204.185 92.320 204.515 ;
        RECT 92.490 204.185 93.370 204.515 ;
        RECT 91.210 204.015 91.455 204.055 ;
        RECT 92.120 204.015 92.320 204.185 ;
        RECT 91.210 203.930 91.610 204.015 ;
        RECT 90.840 203.535 91.090 203.805 ;
        RECT 91.280 203.495 91.610 203.930 ;
        RECT 92.120 203.490 92.450 204.015 ;
        RECT 93.200 203.725 93.370 204.185 ;
        RECT 93.540 204.225 93.860 205.185 ;
        RECT 94.030 204.435 94.220 205.155 ;
        RECT 94.390 204.255 94.560 205.325 ;
        RECT 95.070 205.380 96.175 205.550 ;
        RECT 95.070 204.765 95.240 205.380 ;
        RECT 96.385 205.230 96.635 205.655 ;
        RECT 95.410 204.845 95.940 205.210 ;
        RECT 96.385 205.100 96.690 205.230 ;
        RECT 94.730 204.675 95.240 204.765 ;
        RECT 94.730 204.505 95.600 204.675 ;
        RECT 94.730 204.435 94.900 204.505 ;
        RECT 95.020 204.255 95.220 204.285 ;
        RECT 93.540 203.895 94.005 204.225 ;
        RECT 94.390 203.955 95.220 204.255 ;
        RECT 94.390 203.725 94.560 203.955 ;
        RECT 93.200 203.555 93.985 203.725 ;
        RECT 94.155 203.555 94.560 203.725 ;
        RECT 95.430 203.725 95.600 204.505 ;
        RECT 95.770 204.145 95.940 204.845 ;
        RECT 96.110 204.315 96.350 204.910 ;
        RECT 95.770 203.925 96.295 204.145 ;
        RECT 96.520 203.995 96.690 205.100 ;
        RECT 96.465 203.865 96.690 203.995 ;
        RECT 96.860 203.905 97.140 204.855 ;
        RECT 96.465 203.725 96.635 203.865 ;
        RECT 95.430 203.555 96.105 203.725 ;
        RECT 96.300 203.555 96.635 203.725 ;
        RECT 97.310 203.535 97.495 205.655 ;
        RECT 98.165 205.155 98.335 205.655 ;
        RECT 97.670 204.985 98.335 205.155 ;
        RECT 97.670 203.995 97.900 204.985 ;
        RECT 98.770 204.820 99.105 205.655 ;
        RECT 98.380 204.815 99.105 204.820 ;
        RECT 98.070 204.670 99.105 204.815 ;
        RECT 99.680 204.905 100.010 205.635 ;
        RECT 98.070 204.540 99.005 204.670 ;
        RECT 98.070 204.165 98.420 204.540 ;
        RECT 98.770 204.330 99.005 204.540 ;
        RECT 99.680 204.515 99.950 204.905 ;
        RECT 100.200 204.765 100.530 205.610 ;
        RECT 98.760 204.100 99.005 204.330 ;
        RECT 99.175 204.185 99.950 204.515 ;
        RECT 97.670 203.825 98.335 203.995 ;
        RECT 98.760 203.990 99.025 204.100 ;
        RECT 98.165 203.535 98.335 203.825 ;
        RECT 98.770 203.445 99.025 203.990 ;
        RECT 99.750 203.805 99.950 204.185 ;
        RECT 100.120 204.685 100.530 204.765 ;
        RECT 101.040 205.095 101.380 205.655 ;
        RECT 102.110 205.355 102.995 205.525 ;
        RECT 101.040 204.720 101.940 205.095 ;
        RECT 100.120 204.635 100.355 204.685 ;
        RECT 100.120 204.055 100.310 204.635 ;
        RECT 101.040 204.515 101.230 204.720 ;
        RECT 102.110 204.515 102.280 205.355 ;
        RECT 103.220 205.325 103.470 205.655 ;
        RECT 100.480 204.185 101.230 204.515 ;
        RECT 101.400 204.185 102.280 204.515 ;
        RECT 100.120 204.015 100.365 204.055 ;
        RECT 101.030 204.015 101.230 204.185 ;
        RECT 100.120 203.930 100.520 204.015 ;
        RECT 99.750 203.535 100.000 203.805 ;
        RECT 100.190 203.495 100.520 203.930 ;
        RECT 101.030 203.490 101.360 204.015 ;
        RECT 102.110 203.725 102.280 204.185 ;
        RECT 102.450 204.225 102.770 205.185 ;
        RECT 102.940 204.435 103.130 205.155 ;
        RECT 103.300 204.255 103.470 205.325 ;
        RECT 103.980 205.380 105.085 205.550 ;
        RECT 103.980 204.765 104.150 205.380 ;
        RECT 105.295 205.230 105.545 205.655 ;
        RECT 104.320 204.845 104.850 205.210 ;
        RECT 105.295 205.100 105.600 205.230 ;
        RECT 103.640 204.675 104.150 204.765 ;
        RECT 103.640 204.505 104.510 204.675 ;
        RECT 103.640 204.435 103.810 204.505 ;
        RECT 103.930 204.255 104.130 204.285 ;
        RECT 102.450 203.895 102.915 204.225 ;
        RECT 103.300 203.955 104.130 204.255 ;
        RECT 103.300 203.725 103.470 203.955 ;
        RECT 102.110 203.555 102.895 203.725 ;
        RECT 103.065 203.555 103.470 203.725 ;
        RECT 104.340 203.725 104.510 204.505 ;
        RECT 104.680 204.145 104.850 204.845 ;
        RECT 105.020 204.315 105.260 204.910 ;
        RECT 104.680 203.925 105.205 204.145 ;
        RECT 105.430 203.995 105.600 205.100 ;
        RECT 105.375 203.865 105.600 203.995 ;
        RECT 105.770 203.905 106.050 204.855 ;
        RECT 105.375 203.725 105.545 203.865 ;
        RECT 104.340 203.555 105.015 203.725 ;
        RECT 105.210 203.555 105.545 203.725 ;
        RECT 106.220 203.535 106.405 205.655 ;
        RECT 107.075 205.155 107.245 205.655 ;
        RECT 106.580 204.985 107.245 205.155 ;
        RECT 106.580 203.995 106.810 204.985 ;
        RECT 106.980 204.790 107.330 204.815 ;
        RECT 107.680 204.790 108.015 205.655 ;
        RECT 106.980 204.670 108.015 204.790 ;
        RECT 108.590 204.905 108.920 205.635 ;
        RECT 106.980 204.460 107.915 204.670 ;
        RECT 108.590 204.515 108.860 204.905 ;
        RECT 109.110 204.765 109.440 205.610 ;
        RECT 106.980 204.165 107.330 204.460 ;
        RECT 107.680 204.100 107.915 204.460 ;
        RECT 108.085 204.185 108.860 204.515 ;
        RECT 106.580 203.825 107.245 203.995 ;
        RECT 107.075 203.535 107.245 203.825 ;
        RECT 107.680 203.445 107.935 204.100 ;
        RECT 108.660 203.805 108.860 204.185 ;
        RECT 109.030 204.685 109.440 204.765 ;
        RECT 109.950 205.095 110.290 205.655 ;
        RECT 111.020 205.355 111.905 205.525 ;
        RECT 109.950 204.720 110.850 205.095 ;
        RECT 109.030 204.635 109.265 204.685 ;
        RECT 109.030 204.055 109.220 204.635 ;
        RECT 109.950 204.515 110.140 204.720 ;
        RECT 111.020 204.515 111.190 205.355 ;
        RECT 112.130 205.325 112.380 205.655 ;
        RECT 109.390 204.185 110.140 204.515 ;
        RECT 110.310 204.185 111.190 204.515 ;
        RECT 109.030 204.015 109.275 204.055 ;
        RECT 109.940 204.015 110.140 204.185 ;
        RECT 109.030 203.930 109.430 204.015 ;
        RECT 108.660 203.535 108.910 203.805 ;
        RECT 109.100 203.495 109.430 203.930 ;
        RECT 109.940 203.490 110.270 204.015 ;
        RECT 111.020 203.725 111.190 204.185 ;
        RECT 111.360 204.225 111.680 205.185 ;
        RECT 111.850 204.435 112.040 205.155 ;
        RECT 112.210 204.255 112.380 205.325 ;
        RECT 112.890 205.380 113.995 205.550 ;
        RECT 112.890 204.765 113.060 205.380 ;
        RECT 114.205 205.230 114.455 205.655 ;
        RECT 113.230 204.845 113.760 205.210 ;
        RECT 114.205 205.100 114.510 205.230 ;
        RECT 112.550 204.675 113.060 204.765 ;
        RECT 112.550 204.505 113.420 204.675 ;
        RECT 112.550 204.435 112.720 204.505 ;
        RECT 112.840 204.255 113.040 204.285 ;
        RECT 111.360 203.895 111.825 204.225 ;
        RECT 112.210 203.955 113.040 204.255 ;
        RECT 112.210 203.725 112.380 203.955 ;
        RECT 111.020 203.555 111.805 203.725 ;
        RECT 111.975 203.555 112.380 203.725 ;
        RECT 113.250 203.725 113.420 204.505 ;
        RECT 113.590 204.145 113.760 204.845 ;
        RECT 113.930 204.315 114.170 204.910 ;
        RECT 113.590 203.925 114.115 204.145 ;
        RECT 114.340 203.995 114.510 205.100 ;
        RECT 114.285 203.865 114.510 203.995 ;
        RECT 114.680 203.905 114.960 204.855 ;
        RECT 114.285 203.725 114.455 203.865 ;
        RECT 113.250 203.555 113.925 203.725 ;
        RECT 114.120 203.555 114.455 203.725 ;
        RECT 115.130 203.535 115.315 205.655 ;
        RECT 115.985 205.155 116.155 205.655 ;
        RECT 134.770 205.465 134.980 209.830 ;
        RECT 115.490 204.985 116.155 205.155 ;
        RECT 133.605 205.250 135.805 205.465 ;
        RECT 133.605 205.130 134.575 205.250 ;
        RECT 135.185 205.210 135.805 205.250 ;
        RECT 115.490 203.995 115.720 204.985 ;
        RECT 134.745 204.555 135.075 205.080 ;
        RECT 133.625 204.485 135.075 204.555 ;
        RECT 133.625 204.285 135.725 204.485 ;
        RECT 133.625 204.225 134.355 204.285 ;
        RECT 135.455 204.225 135.725 204.285 ;
        RECT 115.490 203.825 116.155 203.995 ;
        RECT 115.985 203.535 116.155 203.825 ;
        RECT 134.745 202.710 135.075 203.260 ;
        RECT 134.745 202.700 135.770 202.710 ;
        RECT 133.605 202.510 135.770 202.700 ;
        RECT 133.605 202.360 134.540 202.510 ;
        RECT 135.245 202.380 135.770 202.510 ;
        RECT 11.315 201.625 11.485 202.125 ;
        RECT 11.315 201.455 11.980 201.625 ;
        RECT 11.750 200.465 11.980 201.455 ;
        RECT 11.315 200.295 11.980 200.465 ;
        RECT 11.315 200.005 11.485 200.295 ;
        RECT 12.155 200.005 12.340 202.125 ;
        RECT 13.015 201.700 13.265 202.125 ;
        RECT 13.475 201.850 14.580 202.020 ;
        RECT 12.960 201.570 13.265 201.700 ;
        RECT 12.510 200.375 12.790 201.325 ;
        RECT 12.960 200.465 13.130 201.570 ;
        RECT 13.300 200.785 13.540 201.380 ;
        RECT 13.710 201.315 14.240 201.680 ;
        RECT 13.710 200.615 13.880 201.315 ;
        RECT 14.410 201.235 14.580 201.850 ;
        RECT 15.090 201.795 15.340 202.125 ;
        RECT 15.565 201.825 16.450 201.995 ;
        RECT 14.410 201.145 14.920 201.235 ;
        RECT 12.960 200.335 13.185 200.465 ;
        RECT 13.355 200.395 13.880 200.615 ;
        RECT 14.050 200.975 14.920 201.145 ;
        RECT 13.015 200.195 13.185 200.335 ;
        RECT 14.050 200.195 14.220 200.975 ;
        RECT 14.750 200.905 14.920 200.975 ;
        RECT 14.430 200.725 14.630 200.755 ;
        RECT 15.090 200.725 15.260 201.795 ;
        RECT 15.430 200.905 15.620 201.625 ;
        RECT 14.430 200.425 15.260 200.725 ;
        RECT 15.790 200.695 16.110 201.655 ;
        RECT 13.015 200.025 13.350 200.195 ;
        RECT 13.545 200.025 14.220 200.195 ;
        RECT 15.090 200.195 15.260 200.425 ;
        RECT 15.645 200.365 16.110 200.695 ;
        RECT 16.280 200.985 16.450 201.825 ;
        RECT 17.180 201.565 17.520 202.125 ;
        RECT 16.620 201.190 17.520 201.565 ;
        RECT 17.330 200.985 17.520 201.190 ;
        RECT 18.030 201.235 18.360 202.080 ;
        RECT 19.045 201.375 19.375 202.105 ;
        RECT 18.030 201.155 18.440 201.235 ;
        RECT 18.205 201.105 18.440 201.155 ;
        RECT 16.280 200.655 17.160 200.985 ;
        RECT 17.330 200.655 18.080 200.985 ;
        RECT 16.280 200.195 16.450 200.655 ;
        RECT 17.330 200.485 17.530 200.655 ;
        RECT 18.250 200.525 18.440 201.105 ;
        RECT 18.195 200.485 18.440 200.525 ;
        RECT 15.090 200.025 15.495 200.195 ;
        RECT 15.665 200.025 16.450 200.195 ;
        RECT 17.200 199.960 17.530 200.485 ;
        RECT 18.040 200.400 18.440 200.485 ;
        RECT 19.105 200.985 19.375 201.375 ;
        RECT 19.950 201.155 20.285 202.125 ;
        RECT 23.735 201.625 23.905 202.125 ;
        RECT 23.735 201.455 24.400 201.625 ;
        RECT 19.105 200.655 19.900 200.985 ;
        RECT 18.040 199.965 18.370 200.400 ;
        RECT 19.105 200.275 19.305 200.655 ;
        RECT 20.070 200.545 20.285 201.155 ;
        RECT 23.650 200.635 24.000 201.285 ;
        RECT 19.045 200.005 19.305 200.275 ;
        RECT 20.030 199.925 20.285 200.545 ;
        RECT 24.170 200.465 24.400 201.455 ;
        RECT 23.735 200.295 24.400 200.465 ;
        RECT 23.735 200.005 23.905 200.295 ;
        RECT 24.575 200.005 24.760 202.125 ;
        RECT 25.435 201.700 25.685 202.125 ;
        RECT 25.895 201.850 27.000 202.020 ;
        RECT 25.380 201.570 25.685 201.700 ;
        RECT 24.930 200.375 25.210 201.325 ;
        RECT 25.380 200.465 25.550 201.570 ;
        RECT 25.720 200.785 25.960 201.380 ;
        RECT 26.130 201.315 26.660 201.680 ;
        RECT 26.130 200.615 26.300 201.315 ;
        RECT 26.830 201.235 27.000 201.850 ;
        RECT 27.510 201.795 27.760 202.125 ;
        RECT 27.985 201.825 28.870 201.995 ;
        RECT 26.830 201.145 27.340 201.235 ;
        RECT 25.380 200.335 25.605 200.465 ;
        RECT 25.775 200.395 26.300 200.615 ;
        RECT 26.470 200.975 27.340 201.145 ;
        RECT 25.435 200.195 25.605 200.335 ;
        RECT 26.470 200.195 26.640 200.975 ;
        RECT 27.170 200.905 27.340 200.975 ;
        RECT 26.850 200.725 27.050 200.755 ;
        RECT 27.510 200.725 27.680 201.795 ;
        RECT 27.850 200.905 28.040 201.625 ;
        RECT 26.850 200.425 27.680 200.725 ;
        RECT 28.210 200.695 28.530 201.655 ;
        RECT 25.435 200.025 25.770 200.195 ;
        RECT 25.965 200.025 26.640 200.195 ;
        RECT 27.510 200.195 27.680 200.425 ;
        RECT 28.065 200.365 28.530 200.695 ;
        RECT 28.700 200.985 28.870 201.825 ;
        RECT 29.600 201.565 29.940 202.125 ;
        RECT 29.040 201.190 29.940 201.565 ;
        RECT 31.465 201.375 31.795 202.105 ;
        RECT 29.750 200.985 29.940 201.190 ;
        RECT 31.525 200.985 31.795 201.375 ;
        RECT 32.370 201.155 32.705 202.125 ;
        RECT 36.055 201.605 36.225 202.105 ;
        RECT 36.055 201.435 36.720 201.605 ;
        RECT 28.700 200.655 29.580 200.985 ;
        RECT 29.750 200.655 30.500 200.985 ;
        RECT 31.525 200.655 32.320 200.985 ;
        RECT 28.700 200.195 28.870 200.655 ;
        RECT 29.750 200.485 29.950 200.655 ;
        RECT 27.510 200.025 27.915 200.195 ;
        RECT 28.085 200.025 28.870 200.195 ;
        RECT 29.620 199.960 29.950 200.485 ;
        RECT 31.525 200.275 31.725 200.655 ;
        RECT 32.490 200.545 32.705 201.155 ;
        RECT 35.970 200.615 36.320 201.265 ;
        RECT 31.465 200.005 31.725 200.275 ;
        RECT 32.450 199.925 32.705 200.545 ;
        RECT 36.490 200.445 36.720 201.435 ;
        RECT 36.055 200.275 36.720 200.445 ;
        RECT 36.055 199.985 36.225 200.275 ;
        RECT 36.895 199.985 37.080 202.105 ;
        RECT 37.755 201.680 38.005 202.105 ;
        RECT 38.215 201.830 39.320 202.000 ;
        RECT 37.700 201.550 38.005 201.680 ;
        RECT 37.250 200.355 37.530 201.305 ;
        RECT 37.700 200.445 37.870 201.550 ;
        RECT 38.040 200.765 38.280 201.360 ;
        RECT 38.450 201.295 38.980 201.660 ;
        RECT 38.450 200.595 38.620 201.295 ;
        RECT 39.150 201.215 39.320 201.830 ;
        RECT 39.830 201.775 40.080 202.105 ;
        RECT 40.305 201.805 41.190 201.975 ;
        RECT 39.150 201.125 39.660 201.215 ;
        RECT 37.700 200.315 37.925 200.445 ;
        RECT 38.095 200.375 38.620 200.595 ;
        RECT 38.790 200.955 39.660 201.125 ;
        RECT 37.755 200.175 37.925 200.315 ;
        RECT 38.790 200.175 38.960 200.955 ;
        RECT 39.490 200.885 39.660 200.955 ;
        RECT 39.170 200.705 39.370 200.735 ;
        RECT 39.830 200.705 40.000 201.775 ;
        RECT 40.170 200.885 40.360 201.605 ;
        RECT 39.170 200.405 40.000 200.705 ;
        RECT 40.530 200.675 40.850 201.635 ;
        RECT 37.755 200.005 38.090 200.175 ;
        RECT 38.285 200.005 38.960 200.175 ;
        RECT 39.830 200.175 40.000 200.405 ;
        RECT 40.385 200.345 40.850 200.675 ;
        RECT 41.020 200.965 41.190 201.805 ;
        RECT 41.920 201.545 42.260 202.105 ;
        RECT 41.360 201.170 42.260 201.545 ;
        RECT 43.785 201.355 44.115 202.085 ;
        RECT 42.070 200.965 42.260 201.170 ;
        RECT 43.845 200.965 44.115 201.355 ;
        RECT 44.690 201.135 45.025 202.105 ;
        RECT 134.165 201.800 134.540 202.360 ;
        RECT 134.745 201.630 135.075 202.340 ;
        RECT 41.020 200.635 41.900 200.965 ;
        RECT 42.070 200.635 42.820 200.965 ;
        RECT 43.845 200.635 44.640 200.965 ;
        RECT 41.020 200.175 41.190 200.635 ;
        RECT 42.070 200.465 42.270 200.635 ;
        RECT 39.830 200.005 40.235 200.175 ;
        RECT 40.405 200.005 41.190 200.175 ;
        RECT 41.940 199.940 42.270 200.465 ;
        RECT 43.845 200.255 44.045 200.635 ;
        RECT 44.810 200.525 45.025 201.135 ;
        RECT 133.735 201.460 135.705 201.630 ;
        RECT 133.735 200.745 133.905 201.460 ;
        RECT 134.075 200.970 135.365 201.290 ;
        RECT 135.035 200.825 135.365 200.970 ;
        RECT 135.535 200.845 135.705 201.460 ;
        RECT 134.105 200.610 134.825 200.800 ;
        RECT 43.785 199.985 44.045 200.255 ;
        RECT 44.770 199.905 45.025 200.525 ;
        RECT 133.605 200.440 133.935 200.520 ;
        RECT 135.535 200.440 135.705 200.675 ;
        RECT 133.605 200.270 135.705 200.440 ;
        RECT 134.495 199.930 134.825 200.100 ;
        RECT 134.495 199.760 134.755 199.930 ;
        RECT 135.005 199.810 135.305 200.270 ;
        RECT 133.710 199.590 134.755 199.760 ;
        RECT 134.975 199.610 135.305 199.810 ;
        RECT 133.710 198.655 133.880 199.590 ;
        RECT 134.050 199.060 134.415 199.420 ;
        RECT 134.585 199.400 134.755 199.590 ;
        RECT 134.585 199.230 135.705 199.400 ;
        RECT 134.050 198.890 135.335 199.060 ;
        RECT 134.350 198.480 134.945 198.720 ;
        RECT 135.115 198.535 135.335 198.890 ;
        RECT 135.535 198.725 135.705 199.230 ;
        RECT 133.605 198.310 134.160 198.445 ;
        RECT 135.535 198.365 135.705 198.530 ;
        RECT 135.265 198.310 135.705 198.365 ;
        RECT 133.605 198.195 135.705 198.310 ;
        RECT 134.030 198.140 135.395 198.195 ;
        RECT 134.405 197.690 135.355 197.970 ;
        RECT 133.605 197.335 135.725 197.520 ;
        RECT 134.105 196.930 135.435 197.160 ;
        RECT 134.105 196.665 134.275 196.930 ;
        RECT 133.605 196.495 134.275 196.665 ;
        RECT 134.445 196.410 135.095 196.760 ;
        RECT 135.265 196.665 135.435 196.930 ;
        RECT 135.265 196.495 135.725 196.665 ;
        RECT 97.650 195.820 97.950 196.205 ;
        RECT 97.650 195.275 98.040 195.820 ;
        RECT 99.510 195.775 99.735 196.205 ;
        RECT 100.540 195.825 100.710 196.115 ;
        RECT 98.235 195.605 99.735 195.775 ;
        RECT 97.650 194.565 97.820 195.275 ;
        RECT 98.235 195.065 98.405 195.605 ;
        RECT 97.990 194.735 98.405 195.065 ;
        RECT 99.080 195.535 99.735 195.605 ;
        RECT 99.910 195.655 100.710 195.825 ;
        RECT 101.300 195.865 102.170 196.205 ;
        RECT 99.080 194.625 99.250 195.535 ;
        RECT 99.910 195.065 100.080 195.655 ;
        RECT 101.300 195.485 101.470 195.865 ;
        RECT 102.405 195.745 102.575 196.205 ;
        RECT 103.410 195.775 103.580 196.115 ;
        RECT 104.315 195.775 104.485 196.115 ;
        RECT 100.250 195.315 101.470 195.485 ;
        RECT 101.640 195.405 102.100 195.695 ;
        RECT 102.405 195.575 102.965 195.745 ;
        RECT 103.410 195.605 104.485 195.775 ;
        RECT 104.655 195.875 105.335 196.205 ;
        RECT 105.550 195.875 105.800 196.205 ;
        RECT 102.795 195.435 102.965 195.575 ;
        RECT 101.640 195.395 102.605 195.405 ;
        RECT 101.300 195.225 101.470 195.315 ;
        RECT 101.930 195.235 102.605 195.395 ;
        RECT 99.420 195.035 100.080 195.065 ;
        RECT 99.420 194.815 100.255 195.035 ;
        RECT 99.910 194.735 100.255 194.815 ;
        RECT 97.650 194.050 98.030 194.565 ;
        RECT 99.080 194.455 99.735 194.625 ;
        RECT 99.485 194.085 99.735 194.455 ;
        RECT 100.085 194.205 100.255 194.735 ;
        RECT 100.425 194.775 100.965 195.145 ;
        RECT 101.300 195.055 101.705 195.225 ;
        RECT 100.425 194.375 100.665 194.775 ;
        RECT 101.145 194.605 101.365 194.885 ;
        RECT 100.835 194.435 101.365 194.605 ;
        RECT 100.835 194.205 101.005 194.435 ;
        RECT 100.085 194.035 101.005 194.205 ;
        RECT 101.535 194.275 101.705 195.055 ;
        RECT 101.875 194.445 102.225 195.065 ;
        RECT 102.395 194.445 102.605 195.235 ;
        RECT 102.795 195.265 104.295 195.435 ;
        RECT 102.795 194.575 102.965 195.265 ;
        RECT 104.655 195.095 104.825 195.875 ;
        RECT 105.630 195.745 105.800 195.875 ;
        RECT 103.135 194.925 104.825 195.095 ;
        RECT 104.995 195.315 105.460 195.705 ;
        RECT 105.630 195.575 106.025 195.745 ;
        RECT 103.135 194.745 103.305 194.925 ;
        RECT 101.535 193.995 102.485 194.275 ;
        RECT 102.795 194.185 103.055 194.575 ;
        RECT 103.475 194.505 104.265 194.755 ;
        RECT 102.705 194.015 103.055 194.185 ;
        RECT 104.470 194.215 104.640 194.925 ;
        RECT 104.995 194.725 105.165 195.315 ;
        RECT 104.810 194.505 105.165 194.725 ;
        RECT 105.335 194.505 105.685 195.125 ;
        RECT 105.855 194.215 106.025 195.575 ;
        RECT 104.470 194.045 105.325 194.215 ;
        RECT 105.530 194.045 106.025 194.215 ;
        RECT 106.885 194.085 107.055 196.205 ;
        RECT 107.725 195.705 107.980 196.205 ;
        RECT 107.230 195.535 107.980 195.705 ;
        RECT 107.230 194.545 107.460 195.535 ;
        RECT 107.230 194.375 107.980 194.545 ;
        RECT 107.725 194.085 107.980 194.375 ;
        RECT 134.800 192.220 135.010 196.410 ;
        RECT 134.770 192.215 135.020 192.220 ;
        RECT 133.655 192.000 135.855 192.215 ;
        RECT 133.655 191.880 134.625 192.000 ;
        RECT 135.235 191.960 135.855 192.000 ;
        RECT 99.505 191.135 99.805 191.685 ;
        RECT 100.535 191.305 100.985 191.855 ;
        RECT 99.505 190.965 100.445 191.135 ;
        RECT 100.275 190.715 100.445 190.965 ;
        RECT 100.275 190.385 100.565 190.715 ;
        RECT 100.735 190.670 100.985 191.305 ;
        RECT 103.955 191.035 104.285 191.835 ;
        RECT 104.795 191.055 105.125 191.835 ;
        RECT 134.795 191.305 135.125 191.830 ;
        RECT 133.675 191.235 135.125 191.305 ;
        RECT 104.795 191.035 105.560 191.055 ;
        RECT 103.955 190.865 105.560 191.035 ;
        RECT 133.675 191.035 135.775 191.235 ;
        RECT 133.675 190.975 134.405 191.035 ;
        RECT 135.505 190.975 135.775 191.035 ;
        RECT 103.495 190.670 105.125 190.695 ;
        RECT 100.735 190.450 105.125 190.670 ;
        RECT 100.275 190.295 100.445 190.385 ;
        RECT 99.055 190.105 100.445 190.295 ;
        RECT 99.055 189.745 99.385 190.105 ;
        RECT 100.735 189.935 100.985 190.450 ;
        RECT 103.495 190.445 105.125 190.450 ;
        RECT 105.295 190.275 105.560 190.865 ;
        RECT 134.545 190.300 135.380 190.370 ;
        RECT 134.545 190.290 135.815 190.300 ;
        RECT 100.435 189.645 100.985 189.935 ;
        RECT 103.955 190.095 105.560 190.275 ;
        RECT 133.700 190.180 135.815 190.290 ;
        RECT 133.700 190.135 134.675 190.180 ;
        RECT 103.955 189.625 104.285 190.095 ;
        RECT 104.795 189.625 105.125 190.095 ;
        RECT 133.700 189.960 134.625 190.135 ;
        RECT 135.255 190.125 135.815 190.180 ;
        RECT 134.795 189.460 135.125 190.010 ;
        RECT 135.295 189.970 135.815 190.125 ;
        RECT 134.795 189.450 135.820 189.460 ;
        RECT 133.655 189.260 135.820 189.450 ;
        RECT 133.655 189.110 134.590 189.260 ;
        RECT 135.295 189.130 135.820 189.260 ;
        RECT 134.215 188.550 134.590 189.110 ;
        RECT 134.795 188.380 135.125 189.090 ;
        RECT 133.785 188.210 135.755 188.380 ;
        RECT 133.785 187.495 133.955 188.210 ;
        RECT 134.125 187.720 135.415 188.040 ;
        RECT 135.085 187.575 135.415 187.720 ;
        RECT 135.585 187.595 135.755 188.210 ;
        RECT 97.530 187.070 97.830 187.455 ;
        RECT 97.530 186.525 97.920 187.070 ;
        RECT 99.390 187.025 99.615 187.455 ;
        RECT 100.420 187.075 100.590 187.365 ;
        RECT 98.115 186.855 99.615 187.025 ;
        RECT 97.530 185.815 97.700 186.525 ;
        RECT 98.115 186.315 98.285 186.855 ;
        RECT 97.870 185.985 98.285 186.315 ;
        RECT 98.960 186.785 99.615 186.855 ;
        RECT 99.790 186.905 100.590 187.075 ;
        RECT 101.180 187.115 102.050 187.455 ;
        RECT 98.960 185.875 99.130 186.785 ;
        RECT 99.790 186.315 99.960 186.905 ;
        RECT 101.180 186.735 101.350 187.115 ;
        RECT 102.285 186.995 102.455 187.455 ;
        RECT 103.290 187.025 103.460 187.365 ;
        RECT 104.195 187.025 104.365 187.365 ;
        RECT 100.130 186.565 101.350 186.735 ;
        RECT 101.520 186.655 101.980 186.945 ;
        RECT 102.285 186.825 102.845 186.995 ;
        RECT 103.290 186.855 104.365 187.025 ;
        RECT 104.535 187.125 105.215 187.455 ;
        RECT 105.430 187.125 105.680 187.455 ;
        RECT 102.675 186.685 102.845 186.825 ;
        RECT 101.520 186.645 102.485 186.655 ;
        RECT 101.180 186.475 101.350 186.565 ;
        RECT 101.810 186.485 102.485 186.645 ;
        RECT 99.300 186.285 99.960 186.315 ;
        RECT 99.300 186.065 100.135 186.285 ;
        RECT 99.790 185.985 100.135 186.065 ;
        RECT 97.530 185.300 97.910 185.815 ;
        RECT 98.960 185.705 99.615 185.875 ;
        RECT 99.365 185.335 99.615 185.705 ;
        RECT 99.965 185.455 100.135 185.985 ;
        RECT 100.305 186.025 100.845 186.395 ;
        RECT 101.180 186.305 101.585 186.475 ;
        RECT 100.305 185.625 100.545 186.025 ;
        RECT 101.025 185.855 101.245 186.135 ;
        RECT 100.715 185.685 101.245 185.855 ;
        RECT 100.715 185.455 100.885 185.685 ;
        RECT 99.965 185.285 100.885 185.455 ;
        RECT 101.415 185.525 101.585 186.305 ;
        RECT 101.755 185.695 102.105 186.315 ;
        RECT 102.275 185.695 102.485 186.485 ;
        RECT 102.675 186.515 104.175 186.685 ;
        RECT 102.675 185.825 102.845 186.515 ;
        RECT 104.535 186.345 104.705 187.125 ;
        RECT 105.510 186.995 105.680 187.125 ;
        RECT 103.015 186.175 104.705 186.345 ;
        RECT 104.875 186.565 105.340 186.955 ;
        RECT 105.510 186.825 105.905 186.995 ;
        RECT 103.015 185.995 103.185 186.175 ;
        RECT 101.415 185.245 102.365 185.525 ;
        RECT 102.675 185.435 102.935 185.825 ;
        RECT 103.355 185.755 104.145 186.005 ;
        RECT 102.585 185.265 102.935 185.435 ;
        RECT 104.350 185.465 104.520 186.175 ;
        RECT 104.875 185.975 105.045 186.565 ;
        RECT 104.690 185.755 105.045 185.975 ;
        RECT 105.215 185.755 105.565 186.375 ;
        RECT 105.735 185.465 105.905 186.825 ;
        RECT 104.350 185.295 105.205 185.465 ;
        RECT 105.410 185.295 105.905 185.465 ;
        RECT 106.765 185.335 106.935 187.455 ;
        RECT 107.605 186.955 107.860 187.455 ;
        RECT 134.155 187.360 134.875 187.550 ;
        RECT 133.655 187.190 133.985 187.270 ;
        RECT 135.585 187.190 135.755 187.425 ;
        RECT 133.655 187.020 135.755 187.190 ;
        RECT 107.110 186.785 107.860 186.955 ;
        RECT 107.110 185.795 107.340 186.785 ;
        RECT 134.545 186.680 134.875 186.850 ;
        RECT 134.545 186.510 134.805 186.680 ;
        RECT 135.055 186.560 135.355 187.020 ;
        RECT 133.760 186.340 134.805 186.510 ;
        RECT 135.025 186.360 135.355 186.560 ;
        RECT 107.110 185.625 107.860 185.795 ;
        RECT 107.605 185.335 107.860 185.625 ;
        RECT 133.760 185.405 133.930 186.340 ;
        RECT 134.100 185.810 134.465 186.170 ;
        RECT 134.635 186.150 134.805 186.340 ;
        RECT 134.635 185.980 135.755 186.150 ;
        RECT 134.100 185.640 135.385 185.810 ;
        RECT 134.400 185.230 134.995 185.470 ;
        RECT 135.165 185.285 135.385 185.640 ;
        RECT 135.585 185.475 135.755 185.980 ;
        RECT 133.655 185.060 134.210 185.195 ;
        RECT 135.585 185.115 135.755 185.280 ;
        RECT 135.315 185.060 135.755 185.115 ;
        RECT 133.655 184.945 135.755 185.060 ;
        RECT 134.080 184.890 135.445 184.945 ;
        RECT 134.455 184.440 135.405 184.720 ;
        RECT 133.655 184.085 135.775 184.270 ;
        RECT 134.155 183.680 135.485 183.910 ;
        RECT 134.155 183.415 134.325 183.680 ;
        RECT 133.655 183.245 134.325 183.415 ;
        RECT 135.315 183.415 135.485 183.680 ;
        RECT 135.315 183.245 135.775 183.415 ;
        RECT 107.050 27.750 107.850 27.920 ;
        RECT 108.140 27.750 108.940 27.920 ;
        RECT 112.170 27.750 112.970 27.920 ;
        RECT 113.260 27.750 114.060 27.920 ;
        RECT 117.290 27.740 118.090 27.910 ;
        RECT 118.380 27.740 119.180 27.910 ;
        RECT 122.410 27.740 123.210 27.910 ;
        RECT 123.500 27.740 124.300 27.910 ;
        RECT 107.910 24.245 108.080 27.535 ;
        RECT 113.030 24.245 113.200 27.535 ;
        RECT 118.150 24.235 118.320 27.525 ;
        RECT 123.270 24.235 123.440 27.525 ;
        RECT 151.845 27.140 152.175 27.310 ;
        RECT 152.435 27.140 152.765 27.310 ;
        RECT 107.050 23.860 107.850 24.030 ;
        RECT 108.140 23.860 108.940 24.030 ;
        RECT 112.170 23.860 112.970 24.030 ;
        RECT 113.260 23.860 114.060 24.030 ;
        RECT 117.290 23.850 118.090 24.020 ;
        RECT 118.380 23.850 119.180 24.020 ;
        RECT 122.410 23.850 123.210 24.020 ;
        RECT 123.500 23.850 124.300 24.020 ;
        RECT 100.610 21.100 100.940 21.270 ;
        RECT 104.590 21.040 105.340 21.210 ;
        RECT 105.630 21.040 106.380 21.210 ;
        RECT 106.670 21.040 107.420 21.210 ;
        RECT 110.650 21.040 111.400 21.210 ;
        RECT 111.690 21.040 112.440 21.210 ;
        RECT 112.730 21.040 113.480 21.210 ;
        RECT 116.710 21.030 117.460 21.200 ;
        RECT 117.750 21.030 118.500 21.200 ;
        RECT 118.790 21.030 119.540 21.200 ;
        RECT 104.360 18.785 104.530 20.825 ;
        RECT 105.400 18.785 105.570 20.825 ;
        RECT 106.440 18.785 106.610 20.825 ;
        RECT 107.480 18.785 107.650 20.825 ;
        RECT 110.420 18.785 110.590 20.825 ;
        RECT 111.460 18.785 111.630 20.825 ;
        RECT 112.500 18.785 112.670 20.825 ;
        RECT 113.540 18.785 113.710 20.825 ;
        RECT 116.480 18.775 116.650 20.815 ;
        RECT 117.520 18.775 117.690 20.815 ;
        RECT 118.560 18.775 118.730 20.815 ;
        RECT 119.600 18.775 119.770 20.815 ;
        RECT 100.130 18.460 100.460 18.630 ;
        RECT 101.090 18.460 101.420 18.630 ;
        RECT 104.590 18.400 105.340 18.570 ;
        RECT 105.630 18.400 106.380 18.570 ;
        RECT 106.670 18.400 107.420 18.570 ;
        RECT 110.650 18.400 111.400 18.570 ;
        RECT 111.690 18.400 112.440 18.570 ;
        RECT 112.730 18.400 113.480 18.570 ;
        RECT 116.710 18.390 117.460 18.560 ;
        RECT 117.750 18.390 118.500 18.560 ;
        RECT 118.790 18.390 119.540 18.560 ;
        RECT 123.230 18.220 123.400 21.510 ;
        RECT 139.600 20.655 139.770 26.695 ;
        RECT 140.780 20.655 140.950 26.695 ;
        RECT 145.565 26.590 145.895 26.760 ;
        RECT 145.350 20.335 145.520 26.375 ;
        RECT 145.565 19.950 145.895 20.120 ;
        RECT 151.630 19.885 151.800 26.925 ;
        RECT 152.810 19.885 152.980 26.925 ;
        RECT 151.845 19.500 152.175 19.670 ;
        RECT 152.435 19.500 152.765 19.670 ;
        RECT 141.780 17.715 142.110 17.885 ;
        RECT 138.030 17.255 138.360 17.425 ;
        RECT 100.500 16.310 100.830 16.480 ;
        RECT 105.370 16.380 106.120 16.550 ;
        RECT 106.410 16.380 107.160 16.550 ;
        RECT 111.460 16.360 112.210 16.530 ;
        RECT 112.500 16.360 113.250 16.530 ;
        RECT 117.470 16.370 118.220 16.540 ;
        RECT 118.510 16.370 119.260 16.540 ;
        RECT 105.140 13.920 105.310 16.210 ;
        RECT 106.180 13.920 106.350 16.210 ;
        RECT 107.220 13.920 107.390 16.210 ;
        RECT 111.230 13.900 111.400 16.190 ;
        RECT 112.270 13.900 112.440 16.190 ;
        RECT 113.310 13.900 113.480 16.190 ;
        RECT 117.240 13.910 117.410 16.200 ;
        RECT 118.280 13.910 118.450 16.200 ;
        RECT 119.320 13.910 119.490 16.200 ;
        RECT 137.815 15.045 137.985 17.085 ;
        RECT 141.565 15.505 141.735 17.545 ;
        RECT 145.080 15.750 145.580 15.920 ;
        RECT 141.780 15.165 142.110 15.335 ;
        RECT 138.030 14.705 138.360 14.875 ;
        RECT 144.850 14.840 145.020 15.580 ;
        RECT 153.325 15.415 153.495 16.455 ;
        RECT 145.080 14.500 145.580 14.670 ;
        RECT 100.980 13.510 101.310 13.680 ;
        RECT 105.370 13.580 106.120 13.750 ;
        RECT 106.410 13.580 107.160 13.750 ;
        RECT 111.460 13.560 112.210 13.730 ;
        RECT 112.500 13.560 113.250 13.730 ;
        RECT 117.470 13.570 118.220 13.740 ;
        RECT 118.510 13.570 119.260 13.740 ;
        RECT 154.620 11.480 154.790 12.520 ;
        RECT 106.190 8.060 106.360 11.350 ;
        RECT 112.290 8.060 112.460 11.350 ;
        RECT 118.370 8.080 118.540 11.370 ;
      LAYER met1 ;
        RECT 70.585 219.730 70.875 219.775 ;
        RECT 73.705 219.730 73.995 219.775 ;
        RECT 75.595 219.730 75.885 219.775 ;
        RECT 70.585 219.590 75.885 219.730 ;
        RECT 70.585 219.545 70.875 219.590 ;
        RECT 73.705 219.545 73.995 219.590 ;
        RECT 75.595 219.545 75.885 219.590 ;
        RECT 65.000 218.820 65.360 219.150 ;
        RECT 67.360 219.120 67.660 219.170 ;
        RECT 67.290 218.810 67.730 219.120 ;
        RECT 69.280 219.070 69.710 219.180 ;
        RECT 69.280 218.900 69.795 219.070 ;
        RECT 67.360 218.760 67.660 218.810 ;
        RECT 69.505 218.755 69.795 218.900 ;
        RECT 70.585 219.050 70.875 219.095 ;
        RECT 74.165 219.050 74.455 219.095 ;
        RECT 76.000 219.050 76.290 219.095 ;
        RECT 70.585 218.910 76.290 219.050 ;
        RECT 70.585 218.865 70.875 218.910 ;
        RECT 74.165 218.865 74.455 218.910 ;
        RECT 76.000 218.865 76.290 218.910 ;
        RECT 69.205 218.710 69.795 218.755 ;
        RECT 72.445 218.710 73.095 218.755 ;
        RECT 69.205 218.570 73.095 218.710 ;
        RECT 69.205 218.525 69.495 218.570 ;
        RECT 72.445 218.525 73.095 218.570 ;
        RECT 134.720 218.640 135.090 218.890 ;
        RECT 134.720 218.360 135.080 218.640 ;
        RECT 68.610 215.980 68.920 216.020 ;
        RECT 63.830 215.530 64.270 215.840 ;
        RECT 64.530 215.530 64.970 215.840 ;
        RECT 65.760 215.520 66.830 215.780 ;
        RECT 68.610 215.480 69.290 215.980 ;
        RECT 134.780 215.840 135.100 216.330 ;
        RECT 68.610 215.430 68.920 215.480 ;
        RECT 17.200 214.780 17.760 214.810 ;
        RECT 18.190 214.780 18.690 214.850 ;
        RECT 17.200 214.540 18.690 214.780 ;
        RECT 17.200 214.500 17.760 214.540 ;
        RECT 18.190 214.440 18.690 214.540 ;
        RECT 134.445 214.415 134.675 214.705 ;
        RECT 134.105 213.980 134.335 214.270 ;
        RECT 17.300 213.530 17.600 213.540 ;
        RECT 17.270 213.160 17.690 213.530 ;
        RECT 70.585 213.050 70.875 213.095 ;
        RECT 73.705 213.050 73.995 213.095 ;
        RECT 75.595 213.050 75.885 213.095 ;
        RECT 18.860 212.910 19.030 212.920 ;
        RECT 11.800 212.880 12.160 212.900 ;
        RECT 11.790 212.870 12.160 212.880 ;
        RECT 18.540 212.870 19.030 212.910 ;
        RECT 11.790 212.840 19.030 212.870 ;
        RECT 23.310 212.840 23.630 212.940 ;
        RECT 24.590 212.930 24.970 212.970 ;
        RECT 11.790 212.690 23.630 212.840 ;
        RECT 11.790 212.630 12.160 212.690 ;
        RECT 18.540 212.640 23.630 212.690 ;
        RECT 24.570 212.920 24.970 212.930 ;
        RECT 30.890 212.920 31.870 212.970 ;
        RECT 36.500 212.950 36.950 212.990 ;
        RECT 42.810 212.960 43.230 213.030 ;
        RECT 42.810 212.950 43.750 212.960 ;
        RECT 24.570 212.890 31.870 212.920 ;
        RECT 35.150 212.890 35.550 212.920 ;
        RECT 24.570 212.690 35.550 212.890 ;
        RECT 24.570 212.650 24.970 212.690 ;
        RECT 11.800 212.620 12.160 212.630 ;
        RECT 11.385 212.480 11.675 212.525 ;
        RECT 12.575 212.480 12.865 212.525 ;
        RECT 15.095 212.480 15.385 212.525 ;
        RECT 18.860 212.480 19.030 212.640 ;
        RECT 23.310 212.540 23.630 212.640 ;
        RECT 24.590 212.630 24.970 212.650 ;
        RECT 30.890 212.620 35.550 212.690 ;
        RECT 36.500 212.730 43.750 212.950 ;
        RECT 70.585 212.910 75.885 213.050 ;
        RECT 70.585 212.865 70.875 212.910 ;
        RECT 73.705 212.865 73.995 212.910 ;
        RECT 75.595 212.865 75.885 212.910 ;
        RECT 36.500 212.640 36.950 212.730 ;
        RECT 42.810 212.710 43.750 212.730 ;
        RECT 42.810 212.660 43.230 212.710 ;
        RECT 31.620 212.560 35.550 212.620 ;
        RECT 24.185 212.490 24.475 212.535 ;
        RECT 25.375 212.490 25.665 212.535 ;
        RECT 27.895 212.490 28.185 212.535 ;
        RECT 11.385 212.340 15.385 212.480 ;
        RECT 11.385 212.295 11.675 212.340 ;
        RECT 12.575 212.295 12.865 212.340 ;
        RECT 15.095 212.295 15.385 212.340 ;
        RECT 18.760 212.200 19.110 212.480 ;
        RECT 24.185 212.350 28.185 212.490 ;
        RECT 31.620 212.460 31.900 212.560 ;
        RECT 24.185 212.305 24.475 212.350 ;
        RECT 25.375 212.305 25.665 212.350 ;
        RECT 27.895 212.305 28.185 212.350 ;
        RECT 31.570 212.400 31.900 212.460 ;
        RECT 36.095 212.490 36.385 212.535 ;
        RECT 37.285 212.490 37.575 212.535 ;
        RECT 39.805 212.490 40.095 212.535 ;
        RECT 31.570 212.210 31.890 212.400 ;
        RECT 36.095 212.350 40.095 212.490 ;
        RECT 43.530 212.460 43.750 212.710 ;
        RECT 134.150 212.700 134.290 213.980 ;
        RECT 36.095 212.305 36.385 212.350 ;
        RECT 37.285 212.305 37.575 212.350 ;
        RECT 39.805 212.305 40.095 212.350 ;
        RECT 43.490 212.220 43.800 212.460 ;
        RECT 65.250 212.420 65.480 212.470 ;
        RECT 67.390 212.440 67.620 212.460 ;
        RECT 10.990 212.140 11.280 212.185 ;
        RECT 13.090 212.140 13.380 212.185 ;
        RECT 14.660 212.140 14.950 212.185 ;
        RECT 10.990 212.000 14.950 212.140 ;
        RECT 18.860 212.110 19.030 212.200 ;
        RECT 23.790 212.150 24.080 212.195 ;
        RECT 25.890 212.150 26.180 212.195 ;
        RECT 27.460 212.150 27.750 212.195 ;
        RECT 31.620 212.190 31.860 212.210 ;
        RECT 10.990 211.955 11.280 212.000 ;
        RECT 13.090 211.955 13.380 212.000 ;
        RECT 14.660 211.955 14.950 212.000 ;
        RECT 23.790 212.010 27.750 212.150 ;
        RECT 23.790 211.965 24.080 212.010 ;
        RECT 25.890 211.965 26.180 212.010 ;
        RECT 27.460 211.965 27.750 212.010 ;
        RECT 35.700 212.150 35.990 212.195 ;
        RECT 37.800 212.150 38.090 212.195 ;
        RECT 39.370 212.150 39.660 212.195 ;
        RECT 35.700 212.010 39.660 212.150 ;
        RECT 43.530 212.110 43.750 212.220 ;
        RECT 65.190 212.110 65.550 212.420 ;
        RECT 67.290 212.130 67.730 212.440 ;
        RECT 69.280 212.390 69.710 212.520 ;
        RECT 69.280 212.240 69.795 212.390 ;
        RECT 67.390 212.110 67.620 212.130 ;
        RECT 69.505 212.075 69.795 212.240 ;
        RECT 70.585 212.370 70.875 212.415 ;
        RECT 74.165 212.370 74.455 212.415 ;
        RECT 76.000 212.370 76.290 212.415 ;
        RECT 134.105 212.410 134.335 212.700 ;
        RECT 70.585 212.230 76.290 212.370 ;
        RECT 70.585 212.185 70.875 212.230 ;
        RECT 74.165 212.185 74.455 212.230 ;
        RECT 76.000 212.185 76.290 212.230 ;
        RECT 35.700 211.965 35.990 212.010 ;
        RECT 37.800 211.965 38.090 212.010 ;
        RECT 39.370 211.965 39.660 212.010 ;
        RECT 69.205 212.030 69.795 212.075 ;
        RECT 72.445 212.030 73.095 212.075 ;
        RECT 69.205 211.890 73.095 212.030 ;
        RECT 69.205 211.845 69.495 211.890 ;
        RECT 72.445 211.845 73.095 211.890 ;
        RECT 134.150 210.600 134.290 212.410 ;
        RECT 134.490 212.185 134.630 214.415 ;
        RECT 134.445 211.895 134.675 212.185 ;
        RECT 134.490 210.995 134.630 211.895 ;
        RECT 134.830 211.440 135.080 215.840 ;
        RECT 134.800 211.070 135.090 211.440 ;
        RECT 134.445 210.705 134.675 210.995 ;
        RECT 134.105 210.310 134.335 210.600 ;
        RECT 134.670 205.220 135.040 205.470 ;
        RECT 93.980 205.130 94.270 205.175 ;
        RECT 95.550 205.130 95.840 205.175 ;
        RECT 97.650 205.130 97.940 205.175 ;
        RECT 93.980 204.990 97.940 205.130 ;
        RECT 93.980 204.945 94.270 204.990 ;
        RECT 95.550 204.945 95.840 204.990 ;
        RECT 97.650 204.945 97.940 204.990 ;
        RECT 102.890 205.130 103.180 205.175 ;
        RECT 104.460 205.130 104.750 205.175 ;
        RECT 106.560 205.130 106.850 205.175 ;
        RECT 102.890 204.990 106.850 205.130 ;
        RECT 102.890 204.945 103.180 204.990 ;
        RECT 104.460 204.945 104.750 204.990 ;
        RECT 106.560 204.945 106.850 204.990 ;
        RECT 111.800 205.130 112.090 205.175 ;
        RECT 113.370 205.130 113.660 205.175 ;
        RECT 115.470 205.130 115.760 205.175 ;
        RECT 111.800 204.990 115.760 205.130 ;
        RECT 111.800 204.945 112.090 204.990 ;
        RECT 113.370 204.945 113.660 204.990 ;
        RECT 115.470 204.945 115.760 204.990 ;
        RECT 134.670 204.900 135.030 205.220 ;
        RECT 93.545 204.790 93.835 204.835 ;
        RECT 96.065 204.790 96.355 204.835 ;
        RECT 97.255 204.790 97.545 204.835 ;
        RECT 93.545 204.650 97.545 204.790 ;
        RECT 93.545 204.605 93.835 204.650 ;
        RECT 96.065 204.605 96.355 204.650 ;
        RECT 97.255 204.605 97.545 204.650 ;
        RECT 102.455 204.790 102.745 204.835 ;
        RECT 104.975 204.790 105.265 204.835 ;
        RECT 106.165 204.790 106.455 204.835 ;
        RECT 102.455 204.650 106.455 204.790 ;
        RECT 102.455 204.605 102.745 204.650 ;
        RECT 104.975 204.605 105.265 204.650 ;
        RECT 106.165 204.605 106.455 204.650 ;
        RECT 111.365 204.790 111.655 204.835 ;
        RECT 113.885 204.790 114.175 204.835 ;
        RECT 115.075 204.790 115.365 204.835 ;
        RECT 111.365 204.650 115.365 204.790 ;
        RECT 111.365 204.605 111.655 204.650 ;
        RECT 113.885 204.605 114.175 204.650 ;
        RECT 115.075 204.605 115.365 204.650 ;
        RECT 89.140 203.880 89.430 204.490 ;
        RECT 89.830 204.450 90.120 204.490 ;
        RECT 96.860 204.450 97.150 204.510 ;
        RECT 89.830 204.120 97.150 204.450 ;
        RECT 89.830 204.030 90.120 204.120 ;
        RECT 96.860 204.050 97.150 204.120 ;
        RECT 98.730 204.350 99.020 204.390 ;
        RECT 105.770 204.350 106.060 204.410 ;
        RECT 98.730 204.020 106.060 204.350 ;
        RECT 98.730 203.930 99.020 204.020 ;
        RECT 105.770 203.950 106.060 204.020 ;
        RECT 107.670 204.270 107.920 204.320 ;
        RECT 114.710 204.270 114.960 204.330 ;
        RECT 107.670 203.990 114.960 204.270 ;
        RECT 107.670 203.930 107.920 203.990 ;
        RECT 114.710 203.940 114.960 203.990 ;
        RECT 89.140 203.870 91.590 203.880 ;
        RECT 18.150 202.820 19.150 203.820 ;
        RECT 89.140 203.600 91.630 203.870 ;
        RECT 89.140 203.590 91.590 203.600 ;
        RECT 89.180 203.580 91.590 203.590 ;
        RECT 134.710 202.300 135.030 202.710 ;
        RECT 134.710 202.220 135.070 202.300 ;
        RECT 11.710 201.600 12.000 201.645 ;
        RECT 13.810 201.600 14.100 201.645 ;
        RECT 15.380 201.600 15.670 201.645 ;
        RECT 11.710 201.460 15.670 201.600 ;
        RECT 11.710 201.415 12.000 201.460 ;
        RECT 13.810 201.415 14.100 201.460 ;
        RECT 15.380 201.415 15.670 201.460 ;
        RECT 24.130 201.600 24.420 201.645 ;
        RECT 26.230 201.600 26.520 201.645 ;
        RECT 27.800 201.600 28.090 201.645 ;
        RECT 24.130 201.460 28.090 201.600 ;
        RECT 24.130 201.415 24.420 201.460 ;
        RECT 26.230 201.415 26.520 201.460 ;
        RECT 27.800 201.415 28.090 201.460 ;
        RECT 36.450 201.580 36.740 201.625 ;
        RECT 38.550 201.580 38.840 201.625 ;
        RECT 40.120 201.580 40.410 201.625 ;
        RECT 36.450 201.440 40.410 201.580 ;
        RECT 36.450 201.395 36.740 201.440 ;
        RECT 38.550 201.395 38.840 201.440 ;
        RECT 40.120 201.395 40.410 201.440 ;
        RECT 12.105 201.260 12.395 201.305 ;
        RECT 13.295 201.260 13.585 201.305 ;
        RECT 15.815 201.260 16.105 201.305 ;
        RECT 12.105 201.120 16.105 201.260 ;
        RECT 12.105 201.075 12.395 201.120 ;
        RECT 13.295 201.075 13.585 201.120 ;
        RECT 15.815 201.075 16.105 201.120 ;
        RECT 20.050 200.940 20.280 200.990 ;
        RECT 23.620 200.940 24.010 201.320 ;
        RECT 24.525 201.260 24.815 201.305 ;
        RECT 25.715 201.260 26.005 201.305 ;
        RECT 28.235 201.260 28.525 201.305 ;
        RECT 24.525 201.120 28.525 201.260 ;
        RECT 36.845 201.240 37.135 201.285 ;
        RECT 38.035 201.240 38.325 201.285 ;
        RECT 40.555 201.240 40.845 201.285 ;
        RECT 24.525 201.075 24.815 201.120 ;
        RECT 25.715 201.075 26.005 201.120 ;
        RECT 28.235 201.075 28.525 201.120 ;
        RECT 20.050 200.920 24.010 200.940 ;
        RECT 12.500 200.640 24.010 200.920 ;
        RECT 32.480 200.890 32.710 200.900 ;
        RECT 35.970 200.890 36.330 201.220 ;
        RECT 36.845 201.100 40.845 201.240 ;
        RECT 36.845 201.055 37.135 201.100 ;
        RECT 38.035 201.055 38.325 201.100 ;
        RECT 40.555 201.055 40.845 201.100 ;
        RECT 134.425 200.995 134.655 201.285 ;
        RECT 32.480 200.870 36.330 200.890 ;
        RECT 12.500 200.530 20.280 200.640 ;
        RECT 23.620 200.590 24.010 200.640 ;
        RECT 24.860 200.640 36.330 200.870 ;
        RECT 24.860 200.540 32.710 200.640 ;
        RECT 35.970 200.600 36.330 200.640 ;
        RECT 37.200 200.890 37.570 200.920 ;
        RECT 44.780 200.890 45.050 200.950 ;
        RECT 37.200 200.620 45.050 200.890 ;
        RECT 44.780 200.560 45.050 200.620 ;
        RECT 134.085 200.560 134.315 200.850 ;
        RECT 12.500 200.520 12.770 200.530 ;
        RECT 20.050 200.480 20.280 200.530 ;
        RECT 24.870 200.520 25.270 200.540 ;
        RECT 32.480 200.490 32.710 200.540 ;
        RECT 17.990 200.040 18.850 200.320 ;
        RECT 134.130 199.280 134.270 200.560 ;
        RECT 134.085 198.990 134.315 199.280 ;
        RECT 134.130 197.180 134.270 198.990 ;
        RECT 134.470 198.765 134.610 200.995 ;
        RECT 134.425 198.475 134.655 198.765 ;
        RECT 134.470 197.575 134.610 198.475 ;
        RECT 134.840 198.020 135.070 202.220 ;
        RECT 134.790 197.650 135.080 198.020 ;
        RECT 134.425 197.285 134.655 197.575 ;
        RECT 134.085 196.890 134.315 197.180 ;
        RECT 101.815 195.680 102.105 195.725 ;
        RECT 104.935 195.680 105.225 195.725 ;
        RECT 106.825 195.680 107.115 195.725 ;
        RECT 101.815 195.540 107.115 195.680 ;
        RECT 101.815 195.495 102.105 195.540 ;
        RECT 104.935 195.495 105.225 195.540 ;
        RECT 106.825 195.495 107.115 195.540 ;
        RECT 100.735 194.705 101.025 195.020 ;
        RECT 101.815 195.000 102.105 195.045 ;
        RECT 105.395 195.000 105.685 195.045 ;
        RECT 107.230 195.000 107.520 195.045 ;
        RECT 101.815 194.860 107.520 195.000 ;
        RECT 101.815 194.815 102.105 194.860 ;
        RECT 105.395 194.815 105.685 194.860 ;
        RECT 107.230 194.815 107.520 194.860 ;
        RECT 100.435 194.660 101.025 194.705 ;
        RECT 103.675 194.660 104.325 194.705 ;
        RECT 100.435 194.650 104.325 194.660 ;
        RECT 100.435 194.520 104.340 194.650 ;
        RECT 100.435 194.475 100.725 194.520 ;
        RECT 103.640 194.350 104.340 194.520 ;
        RECT 104.290 193.140 106.750 193.150 ;
        RECT 103.560 192.690 106.750 193.140 ;
        RECT 104.290 192.680 106.750 192.690 ;
        RECT 106.100 191.090 106.750 192.680 ;
        RECT 134.710 192.000 135.080 192.250 ;
        RECT 134.720 191.650 135.080 192.000 ;
        RECT 105.290 190.090 106.750 191.090 ;
        RECT 105.290 190.070 105.570 190.090 ;
        RECT 106.100 188.780 106.750 190.090 ;
        RECT 131.760 190.450 132.760 190.580 ;
        RECT 131.760 189.690 132.880 190.450 ;
        RECT 133.900 190.310 134.210 190.410 ;
        RECT 133.900 189.940 135.720 190.310 ;
        RECT 133.900 189.910 135.460 189.940 ;
        RECT 133.900 189.780 134.210 189.910 ;
        RECT 131.760 189.580 132.760 189.690 ;
        RECT 104.240 188.770 106.750 188.780 ;
        RECT 103.520 188.340 106.750 188.770 ;
        RECT 134.850 188.930 135.170 189.420 ;
        RECT 103.520 188.320 104.310 188.340 ;
        RECT 134.475 187.745 134.705 188.035 ;
        RECT 134.135 187.310 134.365 187.600 ;
        RECT 101.695 186.930 101.985 186.975 ;
        RECT 104.815 186.930 105.105 186.975 ;
        RECT 106.705 186.930 106.995 186.975 ;
        RECT 101.695 186.790 106.995 186.930 ;
        RECT 101.695 186.745 101.985 186.790 ;
        RECT 104.815 186.745 105.105 186.790 ;
        RECT 106.705 186.745 106.995 186.790 ;
        RECT 100.615 185.955 100.905 186.270 ;
        RECT 101.695 186.250 101.985 186.295 ;
        RECT 105.275 186.250 105.565 186.295 ;
        RECT 107.110 186.250 107.400 186.295 ;
        RECT 101.695 186.110 107.400 186.250 ;
        RECT 101.695 186.065 101.985 186.110 ;
        RECT 105.275 186.065 105.565 186.110 ;
        RECT 107.110 186.065 107.400 186.110 ;
        RECT 134.180 186.030 134.320 187.310 ;
        RECT 103.610 185.955 104.290 185.960 ;
        RECT 100.315 185.910 100.905 185.955 ;
        RECT 103.555 185.910 104.290 185.955 ;
        RECT 100.315 185.770 104.290 185.910 ;
        RECT 100.315 185.725 100.605 185.770 ;
        RECT 103.555 185.725 104.290 185.770 ;
        RECT 134.135 185.740 134.365 186.030 ;
        RECT 103.610 185.670 104.290 185.725 ;
        RECT 134.180 183.930 134.320 185.740 ;
        RECT 134.520 185.515 134.660 187.745 ;
        RECT 134.475 185.225 134.705 185.515 ;
        RECT 134.520 184.325 134.660 185.225 ;
        RECT 134.850 184.650 135.160 188.930 ;
        RECT 134.860 184.400 135.150 184.650 ;
        RECT 134.475 184.035 134.705 184.325 ;
        RECT 134.135 183.640 134.365 183.930 ;
        RECT 125.260 28.040 125.620 28.050 ;
        RECT 107.080 27.950 125.620 28.040 ;
        RECT 107.070 27.720 125.620 27.950 ;
        RECT 107.080 27.670 125.620 27.720 ;
        RECT 107.880 24.870 108.110 27.515 ;
        RECT 113.000 24.940 113.230 27.515 ;
        RECT 118.120 25.070 118.350 27.505 ;
        RECT 123.220 26.890 123.500 27.670 ;
        RECT 107.800 24.320 108.190 24.870 ;
        RECT 107.880 24.265 108.110 24.320 ;
        RECT 112.920 24.310 113.300 24.940 ;
        RECT 113.000 24.265 113.230 24.310 ;
        RECT 118.030 24.280 118.430 25.070 ;
        RECT 123.240 24.970 123.470 26.890 ;
        RECT 118.120 24.255 118.350 24.280 ;
        RECT 123.160 24.270 123.550 24.970 ;
        RECT 123.240 24.255 123.470 24.270 ;
        RECT 125.260 24.110 125.620 27.670 ;
        RECT 151.865 27.330 152.155 27.340 ;
        RECT 152.455 27.330 152.745 27.340 ;
        RECT 150.670 27.310 152.745 27.330 ;
        RECT 150.670 27.140 153.130 27.310 ;
        RECT 146.940 26.820 147.340 26.850 ;
        RECT 107.050 23.740 125.620 24.110 ;
        RECT 125.260 23.730 125.620 23.740 ;
        RECT 102.180 22.510 102.510 22.530 ;
        RECT 120.020 22.520 120.890 22.540 ;
        RECT 114.680 22.510 120.890 22.520 ;
        RECT 102.180 22.500 103.080 22.510 ;
        RECT 108.790 22.500 120.890 22.510 ;
        RECT 102.180 22.200 120.890 22.500 ;
        RECT 139.570 22.400 139.800 26.675 ;
        RECT 102.180 22.190 120.210 22.200 ;
        RECT 102.180 21.340 102.510 22.190 ;
        RECT 103.040 22.180 120.210 22.190 ;
        RECT 103.040 22.170 114.680 22.180 ;
        RECT 103.040 22.150 108.830 22.170 ;
        RECT 100.620 21.330 102.510 21.340 ;
        RECT 100.620 21.040 102.520 21.330 ;
        RECT 104.620 21.260 108.460 21.270 ;
        RECT 120.530 21.260 120.870 22.200 ;
        RECT 123.200 21.470 123.430 21.490 ;
        RECT 104.620 21.240 108.790 21.260 ;
        RECT 110.680 21.240 114.850 21.260 ;
        RECT 102.180 19.100 102.520 21.040 ;
        RECT 104.610 21.010 108.790 21.240 ;
        RECT 110.670 21.010 114.850 21.240 ;
        RECT 104.620 21.000 108.790 21.010 ;
        RECT 104.330 19.230 104.560 20.805 ;
        RECT 105.270 20.390 105.690 20.820 ;
        RECT 102.180 18.700 102.530 19.100 ;
        RECT 104.220 18.790 104.620 19.230 ;
        RECT 105.370 18.805 105.600 20.390 ;
        RECT 106.410 19.260 106.640 20.805 ;
        RECT 107.450 20.790 107.680 20.805 ;
        RECT 107.370 20.360 107.790 20.790 ;
        RECT 106.340 18.820 106.740 19.260 ;
        RECT 106.410 18.805 106.640 18.820 ;
        RECT 107.450 18.805 107.680 20.360 ;
        RECT 100.160 18.660 102.530 18.700 ;
        RECT 100.150 18.430 102.530 18.660 ;
        RECT 108.460 18.610 108.790 21.000 ;
        RECT 110.680 20.990 114.850 21.010 ;
        RECT 116.700 20.990 120.870 21.260 ;
        RECT 110.390 19.290 110.620 20.805 ;
        RECT 111.370 20.400 111.740 20.810 ;
        RECT 110.310 18.830 110.690 19.290 ;
        RECT 110.390 18.805 110.620 18.830 ;
        RECT 111.430 18.805 111.660 20.400 ;
        RECT 112.470 19.250 112.700 20.805 ;
        RECT 113.510 20.800 113.740 20.805 ;
        RECT 113.440 20.390 113.810 20.800 ;
        RECT 112.390 18.790 112.770 19.250 ;
        RECT 113.510 18.805 113.740 20.390 ;
        RECT 104.620 18.600 108.790 18.610 ;
        RECT 114.520 18.600 114.850 20.990 ;
        RECT 120.530 20.910 120.870 20.990 ;
        RECT 116.450 19.310 116.680 20.795 ;
        RECT 117.490 20.790 117.720 20.795 ;
        RECT 117.440 20.250 117.800 20.790 ;
        RECT 116.370 18.810 116.730 19.310 ;
        RECT 116.450 18.795 116.680 18.810 ;
        RECT 117.490 18.795 117.720 20.250 ;
        RECT 118.530 19.310 118.760 20.795 ;
        RECT 119.570 20.760 119.800 20.795 ;
        RECT 119.500 20.220 119.860 20.760 ;
        RECT 118.450 18.810 118.810 19.310 ;
        RECT 118.530 18.795 118.760 18.810 ;
        RECT 119.570 18.795 119.800 20.220 ;
        RECT 120.540 18.600 120.870 20.910 ;
        RECT 123.140 20.900 123.500 21.470 ;
        RECT 139.400 20.920 139.980 22.400 ;
        RECT 140.750 22.370 140.980 26.675 ;
        RECT 145.560 26.520 147.340 26.820 ;
        RECT 100.160 18.400 102.530 18.430 ;
        RECT 102.180 18.380 102.530 18.400 ;
        RECT 102.190 17.680 102.530 18.380 ;
        RECT 104.610 18.370 108.790 18.600 ;
        RECT 110.670 18.370 114.850 18.600 ;
        RECT 104.620 18.340 108.790 18.370 ;
        RECT 102.150 17.300 102.580 17.680 ;
        RECT 108.460 17.620 108.790 18.340 ;
        RECT 110.680 18.330 114.850 18.370 ;
        RECT 116.700 18.330 120.870 18.600 ;
        RECT 114.520 17.660 114.850 18.330 ;
        RECT 108.460 17.610 112.500 17.620 ;
        RECT 108.460 17.340 112.560 17.610 ;
        RECT 114.480 17.360 114.920 17.660 ;
        RECT 102.190 16.540 102.530 17.300 ;
        RECT 108.460 16.620 108.790 17.340 ;
        RECT 112.140 17.330 112.560 17.340 ;
        RECT 105.400 16.580 108.790 16.620 ;
        RECT 114.520 16.610 114.850 17.360 ;
        RECT 120.540 16.610 120.870 18.330 ;
        RECT 123.200 18.240 123.430 20.900 ;
        RECT 139.570 20.675 139.800 20.920 ;
        RECT 140.620 20.890 141.200 22.370 ;
        RECT 145.320 21.350 145.550 26.355 ;
        RECT 146.940 26.120 147.340 26.520 ;
        RECT 150.670 26.120 151.030 27.140 ;
        RECT 151.865 27.110 152.155 27.140 ;
        RECT 152.455 27.110 152.745 27.140 ;
        RECT 146.940 24.490 147.290 26.120 ;
        RECT 150.680 24.490 151.030 26.120 ;
        RECT 146.940 21.560 151.030 24.490 ;
        RECT 146.940 21.430 147.350 21.560 ;
        RECT 140.750 20.675 140.980 20.890 ;
        RECT 144.420 20.640 145.560 21.350 ;
        RECT 144.420 20.355 145.550 20.640 ;
        RECT 141.580 19.190 142.350 19.290 ;
        RECT 144.420 19.210 145.350 20.355 ;
        RECT 146.940 20.170 147.320 21.430 ;
        RECT 145.590 20.150 147.320 20.170 ;
        RECT 145.585 19.920 147.320 20.150 ;
        RECT 145.590 19.900 147.320 19.920 ;
        RECT 145.590 19.870 147.210 19.900 ;
        RECT 148.210 19.800 149.750 21.560 ;
        RECT 150.740 19.930 151.030 21.560 ;
        RECT 151.600 21.420 151.830 26.905 ;
        RECT 151.550 20.370 152.020 21.420 ;
        RECT 152.780 21.400 153.010 26.905 ;
        RECT 150.710 19.800 151.030 19.930 ;
        RECT 151.600 19.905 151.830 20.370 ;
        RECT 152.700 20.350 153.170 21.400 ;
        RECT 152.780 19.905 153.010 20.350 ;
        RECT 148.210 19.740 149.770 19.800 ;
        RECT 148.230 19.210 149.770 19.740 ;
        RECT 150.670 19.690 151.030 19.800 ;
        RECT 151.865 19.690 152.155 19.700 ;
        RECT 152.455 19.690 152.745 19.700 ;
        RECT 150.670 19.390 152.860 19.690 ;
        RECT 144.420 19.190 149.770 19.210 ;
        RECT 141.580 18.560 149.770 19.190 ;
        RECT 144.420 18.530 145.350 18.560 ;
        RECT 140.400 18.080 140.860 18.110 ;
        RECT 141.230 18.080 142.410 18.100 ;
        RECT 140.400 18.070 142.410 18.080 ;
        RECT 143.260 18.070 143.540 18.080 ;
        RECT 138.420 17.620 139.260 17.710 ;
        RECT 140.400 17.680 143.540 18.070 ;
        RECT 140.400 17.670 141.230 17.680 ;
        RECT 140.400 17.620 140.860 17.670 ;
        RECT 142.410 17.660 143.540 17.680 ;
        RECT 138.060 17.560 140.860 17.620 ;
        RECT 138.010 17.490 140.860 17.560 ;
        RECT 138.000 17.240 140.860 17.490 ;
        RECT 141.535 17.420 141.765 17.525 ;
        RECT 138.050 17.225 138.340 17.240 ;
        RECT 138.810 17.200 140.860 17.240 ;
        RECT 137.785 16.940 138.015 17.065 ;
        RECT 100.520 16.300 102.530 16.540 ;
        RECT 105.390 16.350 108.790 16.580 ;
        RECT 100.520 16.280 102.030 16.300 ;
        RECT 102.190 13.730 102.530 16.300 ;
        RECT 105.110 14.570 105.340 16.190 ;
        RECT 106.150 16.180 106.380 16.190 ;
        RECT 106.090 15.620 106.450 16.180 ;
        RECT 105.040 14.010 105.400 14.570 ;
        RECT 105.110 13.940 105.340 14.010 ;
        RECT 106.150 13.940 106.380 15.620 ;
        RECT 107.190 14.540 107.420 16.190 ;
        RECT 107.140 13.980 107.500 14.540 ;
        RECT 107.190 13.940 107.420 13.980 ;
        RECT 108.460 13.800 108.790 16.350 ;
        RECT 111.460 16.340 114.850 16.610 ;
        RECT 117.480 16.340 120.870 16.610 ;
        RECT 137.630 16.370 138.120 16.940 ;
        RECT 111.480 16.330 112.190 16.340 ;
        RECT 112.520 16.330 113.230 16.340 ;
        RECT 111.200 14.520 111.430 16.170 ;
        RECT 112.160 15.730 112.550 16.180 ;
        RECT 111.120 13.970 111.510 14.520 ;
        RECT 111.200 13.920 111.430 13.970 ;
        RECT 112.240 13.920 112.470 15.730 ;
        RECT 113.280 14.460 113.510 16.170 ;
        RECT 113.220 13.960 113.590 14.460 ;
        RECT 113.280 13.920 113.510 13.960 ;
        RECT 101.000 13.430 102.530 13.730 ;
        RECT 105.390 13.530 108.790 13.800 ;
        RECT 114.520 13.780 114.850 16.340 ;
        RECT 117.210 14.500 117.440 16.180 ;
        RECT 118.180 15.730 118.550 16.180 ;
        RECT 117.140 14.000 117.510 14.500 ;
        RECT 117.210 13.930 117.440 14.000 ;
        RECT 118.250 13.930 118.480 15.730 ;
        RECT 119.290 14.490 119.520 16.180 ;
        RECT 119.210 13.990 119.580 14.490 ;
        RECT 119.290 13.930 119.520 13.990 ;
        RECT 120.540 13.790 120.870 16.340 ;
        RECT 137.785 15.065 138.015 16.370 ;
        RECT 139.470 15.380 140.860 17.200 ;
        RECT 141.250 16.680 141.960 17.420 ;
        RECT 143.260 17.260 143.540 17.660 ;
        RECT 141.535 15.525 141.765 16.680 ;
        RECT 143.260 16.090 143.960 17.260 ;
        RECT 143.260 15.950 145.530 16.090 ;
        RECT 143.260 15.750 145.560 15.950 ;
        RECT 139.470 15.340 142.090 15.380 ;
        RECT 143.260 15.340 143.960 15.750 ;
        RECT 145.100 15.720 145.560 15.750 ;
        RECT 153.050 15.570 153.840 16.470 ;
        RECT 144.820 15.480 145.050 15.560 ;
        RECT 139.470 14.970 143.960 15.340 ;
        RECT 144.650 15.010 145.160 15.480 ;
        RECT 153.295 15.435 153.525 15.570 ;
        RECT 139.470 14.960 140.860 14.970 ;
        RECT 139.460 14.940 140.860 14.960 ;
        RECT 138.050 14.890 138.340 14.905 ;
        RECT 139.460 14.900 140.570 14.940 ;
        RECT 142.030 14.930 143.960 14.970 ;
        RECT 139.460 14.890 139.600 14.900 ;
        RECT 143.500 14.890 143.960 14.930 ;
        RECT 138.000 14.660 139.600 14.890 ;
        RECT 138.070 14.580 139.600 14.660 ;
        RECT 143.720 14.690 143.960 14.890 ;
        RECT 144.820 14.860 145.050 15.010 ;
        RECT 145.100 14.690 145.560 14.700 ;
        RECT 143.720 14.470 145.560 14.690 ;
        RECT 143.720 14.350 145.550 14.470 ;
        RECT 111.450 13.510 114.850 13.780 ;
        RECT 117.470 13.520 120.870 13.790 ;
        RECT 146.750 14.010 147.610 14.160 ;
        RECT 154.680 14.010 155.340 14.110 ;
        RECT 146.750 13.550 155.340 14.010 ;
        RECT 154.680 12.500 155.340 13.550 ;
        RECT 154.590 11.620 155.340 12.500 ;
        RECT 154.590 11.500 154.820 11.620 ;
        RECT 106.160 11.310 106.390 11.330 ;
        RECT 106.090 10.790 106.470 11.310 ;
        RECT 106.160 8.080 106.390 10.790 ;
        RECT 112.180 10.780 112.590 11.340 ;
        RECT 118.340 11.260 118.570 11.350 ;
        RECT 112.260 8.080 112.490 10.780 ;
        RECT 118.320 10.690 118.710 11.260 ;
        RECT 118.340 8.100 118.570 10.690 ;
      LAYER met2 ;
        RECT 65.010 218.770 67.680 219.210 ;
        RECT 67.340 216.650 67.680 218.770 ;
        RECT 63.880 216.360 67.680 216.650 ;
        RECT 63.880 215.480 64.220 216.360 ;
        RECT 69.330 216.030 69.660 219.230 ;
        RECT 134.670 218.410 135.130 218.690 ;
        RECT 134.770 218.000 135.080 218.410 ;
        RECT 134.760 216.280 135.090 218.000 ;
        RECT 64.580 215.810 64.920 215.890 ;
        RECT 64.580 215.520 67.680 215.810 ;
        RECT 64.580 215.480 64.920 215.520 ;
        RECT 17.250 214.450 17.710 214.860 ;
        RECT 17.310 213.580 17.630 214.450 ;
        RECT 17.310 213.430 17.640 213.580 ;
        RECT 17.320 213.110 17.640 213.430 ;
        RECT 11.850 212.570 12.110 212.950 ;
        RECT 18.590 212.590 18.870 212.960 ;
        RECT 24.640 212.580 24.920 213.020 ;
        RECT 30.940 212.570 31.220 213.020 ;
        RECT 36.550 212.590 36.900 213.040 ;
        RECT 42.860 212.610 43.180 213.080 ;
        RECT 67.340 212.480 67.680 215.520 ;
        RECT 68.660 215.430 69.660 216.030 ;
        RECT 134.730 215.890 135.150 216.280 ;
        RECT 65.210 212.060 67.680 212.480 ;
        RECT 69.330 212.190 69.660 215.430 ;
        RECT 134.620 204.950 135.080 205.230 ;
        RECT 18.430 203.270 18.790 203.310 ;
        RECT 18.420 199.990 18.800 203.270 ;
        RECT 134.710 202.660 135.000 204.950 ;
        RECT 134.660 202.270 135.080 202.660 ;
        RECT 103.620 193.190 104.330 194.740 ;
        RECT 103.610 193.160 104.330 193.190 ;
        RECT 103.610 192.640 104.300 193.160 ;
        RECT 134.670 191.700 135.130 191.980 ;
        RECT 134.730 191.640 135.130 191.700 ;
        RECT 132.840 190.400 133.920 190.410 ;
        RECT 132.420 190.360 133.920 190.400 ;
        RECT 132.420 189.830 134.260 190.360 ;
        RECT 134.790 190.310 135.130 191.640 ;
        RECT 134.730 189.910 135.170 190.310 ;
        RECT 134.730 189.900 135.120 189.910 ;
        RECT 132.420 189.760 133.920 189.830 ;
        RECT 132.420 189.740 132.930 189.760 ;
        RECT 134.790 189.420 135.120 189.900 ;
        RECT 134.790 189.370 135.170 189.420 ;
        RECT 134.790 189.330 135.220 189.370 ;
        RECT 134.800 188.980 135.220 189.330 ;
        RECT 103.570 188.320 104.260 188.820 ;
        RECT 103.570 185.770 104.310 188.320 ;
        RECT 103.580 185.660 104.310 185.770 ;
        RECT 103.660 185.620 104.240 185.660 ;
        RECT 118.080 25.100 118.380 25.120 ;
        RECT 112.970 24.970 113.250 24.990 ;
        RECT 107.850 24.350 108.140 24.920 ;
        RECT 107.850 24.270 108.150 24.350 ;
        RECT 107.860 22.680 108.150 24.270 ;
        RECT 106.680 22.390 108.150 22.680 ;
        RECT 105.320 20.830 105.640 20.870 ;
        RECT 105.320 20.810 105.650 20.830 ;
        RECT 106.680 20.810 107.040 22.390 ;
        RECT 107.860 22.380 108.150 22.390 ;
        RECT 107.420 20.810 107.740 20.840 ;
        RECT 111.420 20.820 111.690 20.860 ;
        RECT 112.940 20.820 113.310 24.970 ;
        RECT 118.080 24.230 118.490 25.100 ;
        RECT 123.210 24.970 123.500 25.020 ;
        RECT 113.490 20.820 113.760 20.850 ;
        RECT 105.320 20.370 107.780 20.810 ;
        RECT 111.420 20.370 113.760 20.820 ;
        RECT 105.320 20.340 105.640 20.370 ;
        RECT 107.420 20.310 107.740 20.370 ;
        RECT 111.420 20.350 111.690 20.370 ;
        RECT 113.490 20.340 113.760 20.370 ;
        RECT 117.490 20.730 117.750 20.840 ;
        RECT 118.100 20.730 118.490 24.230 ;
        RECT 123.170 20.900 123.500 24.970 ;
        RECT 139.450 22.340 139.930 22.450 ;
        RECT 140.670 22.340 141.150 22.420 ;
        RECT 139.450 21.010 141.220 22.340 ;
        RECT 139.050 20.940 141.220 21.010 ;
        RECT 151.600 21.320 151.970 21.470 ;
        RECT 152.750 21.320 153.120 21.450 ;
        RECT 123.190 20.850 123.450 20.900 ;
        RECT 119.550 20.730 119.810 20.810 ;
        RECT 117.490 20.210 119.840 20.730 ;
        RECT 117.490 20.200 117.750 20.210 ;
        RECT 119.550 20.170 119.810 20.210 ;
        RECT 104.270 19.250 104.570 19.280 ;
        RECT 106.390 19.250 106.690 19.310 ;
        RECT 104.270 18.850 106.690 19.250 ;
        RECT 104.270 18.740 104.570 18.850 ;
        RECT 106.090 18.770 106.690 18.850 ;
        RECT 110.360 19.290 110.640 19.340 ;
        RECT 116.420 19.310 116.680 19.360 ;
        RECT 118.500 19.310 118.760 19.360 ;
        RECT 112.440 19.290 112.720 19.300 ;
        RECT 110.360 18.780 112.730 19.290 ;
        RECT 116.420 18.800 118.790 19.310 ;
        RECT 102.200 17.670 102.530 17.730 ;
        RECT 106.090 17.670 106.440 18.770 ;
        RECT 102.200 17.310 106.440 17.670 ;
        RECT 112.200 18.740 112.720 18.780 ;
        RECT 116.420 18.760 116.680 18.800 ;
        RECT 118.180 18.760 118.760 18.800 ;
        RECT 139.050 18.780 140.040 20.940 ;
        RECT 140.670 20.840 141.150 20.940 ;
        RECT 151.600 20.740 153.240 21.320 ;
        RECT 151.600 20.390 153.680 20.740 ;
        RECT 151.600 20.320 151.970 20.390 ;
        RECT 112.200 17.660 112.500 18.740 ;
        RECT 114.530 17.660 114.870 17.710 ;
        RECT 118.180 17.660 118.500 18.760 ;
        RECT 136.940 18.560 140.040 18.780 ;
        RECT 136.930 18.260 140.040 18.560 ;
        RECT 140.860 19.340 142.110 19.360 ;
        RECT 140.860 18.510 142.300 19.340 ;
        RECT 152.500 18.830 153.680 20.390 ;
        RECT 136.930 18.240 139.100 18.260 ;
        RECT 102.200 17.250 102.530 17.310 ;
        RECT 106.090 17.300 106.440 17.310 ;
        RECT 106.100 15.620 106.430 17.300 ;
        RECT 112.190 17.280 112.510 17.660 ;
        RECT 114.520 17.360 118.530 17.660 ;
        RECT 136.930 17.600 137.890 18.240 ;
        RECT 138.060 18.210 139.100 18.240 ;
        RECT 138.520 17.760 139.100 18.210 ;
        RECT 140.860 18.160 142.130 18.510 ;
        RECT 140.860 18.130 141.760 18.160 ;
        RECT 114.530 17.310 114.870 17.360 ;
        RECT 112.200 15.710 112.500 17.280 ;
        RECT 118.180 15.730 118.500 17.360 ;
        RECT 136.930 17.210 137.870 17.600 ;
        RECT 138.470 17.390 139.210 17.760 ;
        RECT 140.860 17.640 141.750 18.130 ;
        RECT 152.520 17.970 153.670 18.830 ;
        RECT 140.860 17.470 141.760 17.640 ;
        RECT 136.930 17.080 137.910 17.210 ;
        RECT 136.930 16.990 138.050 17.080 ;
        RECT 136.930 16.460 138.070 16.990 ;
        RECT 140.860 16.670 141.910 17.470 ;
        RECT 152.520 17.060 153.690 17.970 ;
        RECT 144.800 16.680 145.290 16.690 ;
        RECT 146.360 16.680 147.030 16.710 ;
        RECT 141.300 16.630 141.910 16.670 ;
        RECT 137.410 16.420 138.070 16.460 ;
        RECT 137.680 16.320 138.070 16.420 ;
        RECT 144.780 16.250 147.030 16.680 ;
        RECT 112.210 15.680 112.500 15.710 ;
        RECT 118.230 15.680 118.500 15.730 ;
        RECT 106.140 15.570 106.400 15.620 ;
        RECT 144.800 15.530 145.290 16.250 ;
        RECT 144.700 15.430 145.290 15.530 ;
        RECT 144.700 15.110 145.310 15.430 ;
        RECT 144.700 14.960 145.110 15.110 ;
        RECT 105.090 14.590 105.350 14.620 ;
        RECT 105.090 13.970 107.460 14.590 ;
        RECT 111.170 14.500 111.460 14.570 ;
        RECT 113.270 14.500 113.540 14.510 ;
        RECT 105.090 13.960 105.350 13.970 ;
        RECT 106.120 10.790 106.420 13.970 ;
        RECT 107.190 13.930 107.450 13.970 ;
        RECT 111.170 13.960 113.550 14.500 ;
        RECT 117.190 14.490 117.460 14.550 ;
        RECT 119.260 14.490 119.530 14.540 ;
        RECT 117.190 13.990 119.590 14.490 ;
        RECT 146.360 14.210 147.030 16.250 ;
        RECT 152.490 16.520 153.670 17.060 ;
        RECT 152.490 15.650 153.790 16.520 ;
        RECT 153.100 15.520 153.790 15.650 ;
        RECT 111.170 13.920 111.460 13.960 ;
        RECT 106.140 10.740 106.420 10.790 ;
        RECT 112.210 10.780 112.540 13.960 ;
        RECT 113.270 13.910 113.540 13.960 ;
        RECT 117.190 13.950 117.460 13.990 ;
        RECT 118.350 11.230 118.680 13.990 ;
        RECT 119.260 13.940 119.530 13.990 ;
        RECT 146.360 13.580 147.560 14.210 ;
        RECT 146.800 13.500 147.560 13.580 ;
        RECT 112.230 10.730 112.540 10.780 ;
        RECT 118.370 10.670 118.680 11.230 ;
        RECT 118.370 10.640 118.660 10.670 ;
  END
END tt_um_vks_pll
END LIBRARY

