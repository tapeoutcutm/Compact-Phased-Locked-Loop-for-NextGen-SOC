magic
tech sky130A
magscale 1 2
timestamp 1712737205
<< nwell >>
rect 3772 106 4080 444
rect 2558 -758 2914 -434
rect 3468 -630 3650 -432
rect 3818 -1646 4036 -1300
<< pwell >>
rect 3810 -136 3966 56
rect 3436 -996 3608 -804
rect 3850 -1874 3986 -1708
<< psubdiff >>
rect 3836 -24 3940 30
rect 3836 -58 3867 -24
rect 3901 -58 3940 -24
rect 3836 -110 3940 -58
rect 3462 -884 3582 -830
rect 3462 -918 3504 -884
rect 3538 -918 3582 -884
rect 3462 -970 3582 -918
rect 3876 -1776 3960 -1734
rect 3876 -1810 3900 -1776
rect 3934 -1810 3960 -1776
rect 3876 -1848 3960 -1810
<< nsubdiff >>
rect 3842 298 3922 344
rect 3842 264 3866 298
rect 3900 264 3922 298
rect 3842 220 3922 264
rect 3528 -514 3614 -468
rect 3528 -548 3554 -514
rect 3588 -548 3614 -514
rect 3528 -594 3614 -548
rect 3882 -1464 3968 -1416
rect 3882 -1498 3904 -1464
rect 3938 -1498 3968 -1464
rect 3882 -1550 3968 -1498
<< psubdiffcont >>
rect 3867 -58 3901 -24
rect 3504 -918 3538 -884
rect 3900 -1810 3934 -1776
<< nsubdiffcont >>
rect 3866 264 3900 298
rect 3554 -548 3588 -514
rect 3904 -1498 3938 -1464
<< locali >>
rect 3846 416 3916 420
rect 1886 314 1938 386
rect 3804 380 3916 416
rect 3846 298 3916 380
rect 3846 264 3866 298
rect 3900 264 3916 298
rect 3846 226 3916 264
rect 1108 169 1674 176
rect 1108 63 1129 169
rect 1235 63 1674 169
rect 1108 56 1674 63
rect 3448 111 3498 144
rect 3448 77 3456 111
rect 3490 77 3498 111
rect 3448 44 3498 77
rect 3834 -24 3938 28
rect 3834 -58 3867 -24
rect 3901 -58 3938 -24
rect 3834 -120 3938 -58
rect 3756 -166 3938 -120
rect 3456 -494 3608 -450
rect 3534 -514 3608 -494
rect 3534 -548 3554 -514
rect 3588 -548 3608 -514
rect 3534 -584 3608 -548
rect 2114 -689 2158 -688
rect 2114 -723 2119 -689
rect 2153 -723 2158 -689
rect 2114 -761 2158 -723
rect 3358 -756 3448 -748
rect 3210 -759 3260 -756
rect 2114 -795 2119 -761
rect 2153 -795 2158 -761
rect 2114 -833 2158 -795
rect 2474 -804 3070 -760
rect 3210 -793 3218 -759
rect 3252 -793 3260 -759
rect 3210 -796 3260 -793
rect 3358 -790 3386 -756
rect 3420 -790 3448 -756
rect 3358 -798 3448 -790
rect 2114 -867 2119 -833
rect 2153 -867 2158 -833
rect 2114 -868 2158 -867
rect 3466 -884 3574 -834
rect 3466 -918 3504 -884
rect 3538 -918 3574 -884
rect 3466 -998 3574 -918
rect 3426 -1034 3574 -998
rect 1908 -1438 1960 -1366
rect 3824 -1376 3968 -1330
rect 3882 -1464 3964 -1376
rect 3882 -1498 3904 -1464
rect 3938 -1498 3964 -1464
rect 3882 -1552 3964 -1498
rect 1132 -1582 1704 -1572
rect 1132 -1688 1159 -1582
rect 1265 -1688 1704 -1582
rect 1132 -1698 1704 -1688
rect 1274 -1700 1704 -1698
rect 3472 -1644 3480 -1610
rect 3514 -1644 3522 -1610
rect 3472 -1682 3522 -1644
rect 3472 -1716 3480 -1682
rect 3514 -1716 3522 -1682
rect 3876 -1776 3956 -1736
rect 3876 -1810 3900 -1776
rect 3934 -1810 3956 -1776
rect 3876 -1876 3956 -1810
rect 3766 -1914 3960 -1876
<< viali >>
rect 1129 63 1235 169
rect 3456 77 3490 111
rect 2119 -723 2153 -689
rect 2119 -795 2153 -761
rect 3218 -793 3252 -759
rect 3386 -790 3420 -756
rect 2119 -867 2153 -833
rect 1159 -1688 1265 -1582
rect 3480 -1644 3514 -1610
rect 3480 -1716 3514 -1682
<< metal1 >>
rect 1354 446 1554 646
rect 1354 354 1684 446
rect 1024 182 1224 214
rect 1024 169 1268 182
rect 1024 63 1129 169
rect 1235 63 1268 169
rect 1024 50 1268 63
rect 1024 14 1224 50
rect 1354 -450 1564 354
rect 4156 156 4356 198
rect 3442 111 4356 156
rect 3442 77 3456 111
rect 3490 96 4356 111
rect 3490 77 3551 96
rect 3442 44 3551 77
rect 3603 44 3615 96
rect 3667 44 4356 96
rect 2354 32 2494 36
rect 3442 32 4356 44
rect 2354 -20 2366 32
rect 2418 -20 2430 32
rect 2482 -20 2494 32
rect 3444 28 4356 32
rect 4156 -2 4356 28
rect 2354 -24 2494 -20
rect 3924 -102 4126 -100
rect 3752 -194 4126 -102
rect 3536 -255 3684 -248
rect 1354 -502 1412 -450
rect 1464 -502 1564 -450
rect 1354 -1306 1564 -502
rect 1872 -266 2364 -264
rect 1872 -285 2510 -266
rect 1872 -337 2373 -285
rect 2425 -337 2437 -285
rect 2489 -337 2510 -285
rect 3536 -307 3552 -255
rect 3604 -307 3616 -255
rect 3668 -307 3684 -255
rect 3536 -314 3684 -307
rect 1872 -356 2510 -337
rect 1872 -358 2364 -356
rect 1872 -676 2002 -358
rect 2074 -446 2182 -426
rect 2074 -498 2102 -446
rect 2154 -498 2182 -446
rect 2074 -518 2182 -498
rect 2480 -516 2970 -426
rect 1872 -689 2164 -676
rect 1872 -723 2119 -689
rect 2153 -723 2164 -689
rect 1872 -761 2164 -723
rect 3546 -742 3674 -314
rect 1872 -795 2119 -761
rect 2153 -795 2164 -761
rect 1872 -833 2164 -795
rect 1872 -867 2119 -833
rect 2153 -867 2164 -833
rect 3198 -759 3272 -750
rect 3198 -793 3218 -759
rect 3252 -793 3272 -759
rect 3198 -866 3272 -793
rect 3346 -756 3674 -742
rect 3346 -790 3386 -756
rect 3420 -790 3674 -756
rect 3346 -804 3674 -790
rect 1872 -876 2164 -867
rect 1872 -1138 2002 -876
rect 2108 -880 2164 -876
rect 3188 -867 3284 -866
rect 3188 -919 3210 -867
rect 3262 -919 3284 -867
rect 3188 -920 3284 -919
rect 3924 -966 4126 -194
rect 2468 -1064 4126 -966
rect 1872 -1140 2374 -1138
rect 1872 -1159 2518 -1140
rect 1872 -1211 2381 -1159
rect 2433 -1211 2445 -1159
rect 2497 -1211 2518 -1159
rect 1872 -1226 2518 -1211
rect 2360 -1230 2518 -1226
rect 1354 -1398 1694 -1306
rect 1632 -1400 1694 -1398
rect 1046 -1566 1246 -1534
rect 1046 -1582 1304 -1566
rect 1046 -1688 1159 -1582
rect 1265 -1688 1304 -1582
rect 1046 -1704 1304 -1688
rect 3466 -1600 3528 -1598
rect 3466 -1605 3814 -1600
rect 3466 -1610 3734 -1605
rect 3466 -1644 3480 -1610
rect 3514 -1644 3734 -1610
rect 3466 -1657 3734 -1644
rect 3786 -1657 3814 -1605
rect 3466 -1669 3814 -1657
rect 3466 -1682 3734 -1669
rect 1046 -1734 1246 -1704
rect 2364 -1705 2500 -1702
rect 2364 -1757 2374 -1705
rect 2426 -1757 2438 -1705
rect 2490 -1757 2500 -1705
rect 3466 -1716 3480 -1682
rect 3514 -1716 3734 -1682
rect 3466 -1721 3734 -1716
rect 3786 -1721 3814 -1669
rect 3466 -1726 3814 -1721
rect 3466 -1728 3528 -1726
rect 2364 -1760 2500 -1757
rect 3924 -1850 4126 -1064
rect 4296 -1596 4496 -1570
rect 4254 -1602 4496 -1596
rect 4196 -1607 4496 -1602
rect 4196 -1659 4224 -1607
rect 4276 -1659 4496 -1607
rect 4196 -1671 4496 -1659
rect 4196 -1723 4224 -1671
rect 4276 -1723 4496 -1671
rect 4196 -1728 4496 -1723
rect 4254 -1734 4496 -1728
rect 4296 -1770 4496 -1734
rect 3774 -1942 4126 -1850
rect 3924 -2182 4126 -1942
<< via1 >>
rect 3551 44 3603 96
rect 3615 44 3667 96
rect 2366 -20 2418 32
rect 2430 -20 2482 32
rect 1412 -502 1464 -450
rect 2373 -337 2425 -285
rect 2437 -337 2489 -285
rect 3552 -307 3604 -255
rect 3616 -307 3668 -255
rect 2102 -498 2154 -446
rect 3210 -919 3262 -867
rect 2381 -1211 2433 -1159
rect 2445 -1211 2497 -1159
rect 3734 -1657 3786 -1605
rect 2374 -1757 2426 -1705
rect 2438 -1757 2490 -1705
rect 3734 -1721 3786 -1669
rect 4224 -1659 4276 -1607
rect 4224 -1723 4276 -1671
<< metal2 >>
rect 3546 96 3672 108
rect 2356 32 2498 54
rect 2356 -20 2366 32
rect 2418 -20 2430 32
rect 2482 -20 2498 32
rect 2356 -256 2498 -20
rect 3546 44 3551 96
rect 3603 44 3615 96
rect 3667 44 3672 96
rect 3546 -238 3672 44
rect 3546 -255 3674 -238
rect 2356 -262 2500 -256
rect 2362 -285 2500 -262
rect 2362 -337 2373 -285
rect 2425 -337 2437 -285
rect 2489 -337 2500 -285
rect 3546 -307 3552 -255
rect 3604 -307 3616 -255
rect 3668 -307 3674 -255
rect 3546 -324 3674 -307
rect 2362 -366 2500 -337
rect 1394 -426 1482 -420
rect 2084 -426 2172 -416
rect 1394 -446 2172 -426
rect 1394 -450 2102 -446
rect 1394 -502 1412 -450
rect 1464 -498 2102 -450
rect 2154 -498 2172 -446
rect 1464 -502 2172 -498
rect 1394 -522 2172 -502
rect 1394 -532 1482 -522
rect 2084 -528 2172 -522
rect 3198 -867 3274 -856
rect 3198 -919 3210 -867
rect 3262 -919 3274 -867
rect 3198 -920 3274 -919
rect 2370 -1159 2508 -1130
rect 2370 -1211 2381 -1159
rect 2433 -1211 2445 -1159
rect 2497 -1211 2508 -1159
rect 2370 -1230 2508 -1211
rect 3196 -1154 3274 -920
rect 3196 -1220 3790 -1154
rect 2360 -1705 2508 -1230
rect 2360 -1757 2374 -1705
rect 2426 -1757 2438 -1705
rect 2490 -1740 2508 -1705
rect 3716 -1590 3788 -1220
rect 3716 -1598 3804 -1590
rect 3716 -1602 4030 -1598
rect 4206 -1602 4294 -1592
rect 3716 -1605 4294 -1602
rect 3716 -1657 3734 -1605
rect 3786 -1607 4294 -1605
rect 3786 -1657 4224 -1607
rect 3716 -1659 4224 -1657
rect 4276 -1659 4294 -1607
rect 3716 -1669 4294 -1659
rect 3716 -1721 3734 -1669
rect 3786 -1671 4294 -1669
rect 3786 -1721 4224 -1671
rect 3716 -1723 4224 -1721
rect 4276 -1723 4294 -1671
rect 3716 -1730 4294 -1723
rect 3716 -1732 4030 -1730
rect 3716 -1736 3804 -1732
rect 4206 -1738 4294 -1730
rect 2490 -1757 2506 -1740
rect 2360 -1762 2506 -1757
rect 2374 -1770 2490 -1762
use sky130_fd_sc_hd__dfrbp_2  x1
timestamp 1712737205
transform 1 0 1608 0 1 -146
box -38 -48 2246 592
use sky130_fd_sc_hd__dfrbp_2  x2
timestamp 1712737205
transform 1 0 1632 0 1 -1896
box -38 -48 2246 592
use sky130_fd_sc_hd__and2_2  x3
timestamp 1712737205
transform -1 0 3468 0 1 -1016
box -38 -48 590 592
use sky130_fd_sc_hd__inv_4  x4
timestamp 1712737205
transform -1 0 2544 0 1 -1020
box -38 -48 498 592
<< labels >>
flabel metal1 s 1024 14 1224 214 0 FreeSans 500 0 0 0 A
port 1 nsew
flabel metal1 s 4156 -2 4356 198 0 FreeSans 500 0 0 0 QA
port 2 nsew
flabel metal1 s 1354 446 1554 646 0 FreeSans 500 0 0 0 VDD
port 3 nsew
flabel metal1 s 3926 -2182 4126 -1982 0 FreeSans 500 0 0 0 VSS
port 4 nsew
flabel metal1 s 4296 -1770 4496 -1570 0 FreeSans 500 0 0 0 QB
port 5 nsew
flabel metal1 s 1046 -1734 1246 -1534 0 FreeSans 500 0 0 0 B
port 6 nsew
<< end >>
