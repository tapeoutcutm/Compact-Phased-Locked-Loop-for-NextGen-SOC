magic
tech sky130A
magscale 1 2
timestamp 1709898966
<< error_p >>
rect 17377 2322 17383 2327
rect 17371 2315 17376 2321
rect 17371 2023 17376 2029
rect 17377 2017 17383 2022
<< error_s >>
rect 22866 2732 22886 2958
rect 22894 2760 22914 2930
<< metal1 >>
rect 118 4162 128 5146
rect 600 4859 610 5146
rect 600 4617 25860 4859
rect 600 4162 610 4617
rect 22100 4234 22938 4434
rect 22100 636 22300 4234
rect 26162 4200 31478 4412
rect 22634 2726 22644 3028
rect 22886 2726 22896 3028
rect 26215 2739 27035 2925
rect 23024 2342 23284 2540
rect 22996 2006 23006 2342
rect 23306 2006 23316 2342
rect 26849 959 27035 2739
rect 26849 710 27036 959
rect 22378 636 22388 670
rect 22100 450 22388 636
rect 22300 436 22388 450
rect 22378 428 22388 436
rect 22644 428 22654 670
rect 26804 274 26814 710
rect 27086 274 27096 710
rect 31266 708 31478 4200
rect 31216 358 31226 708
rect 31512 358 31522 708
rect 26849 259 27036 274
rect 26849 251 27035 259
<< via1 >>
rect 128 4162 600 5146
rect 22644 2726 22886 3028
rect 23006 2006 23306 2342
rect 22388 428 22644 670
rect 26814 274 27086 710
rect 31226 358 31512 708
<< metal2 >>
rect 128 5146 600 5156
rect 128 4152 600 4162
rect 18026 3096 18252 3106
rect 22644 3028 22886 3038
rect 18252 2764 22644 2964
rect 18026 2730 18252 2740
rect 22644 2716 22886 2726
rect 23006 2342 23306 2352
rect 23006 1996 23306 2006
rect 26814 710 27086 720
rect 22388 670 22644 680
rect 22388 418 22644 428
rect 31226 708 31512 718
rect 31226 348 31512 358
rect 26814 264 27086 274
<< via2 >>
rect 128 4162 600 5146
rect 18026 2740 18252 3096
rect 23006 2006 23306 2342
rect 22388 428 22644 670
rect 26814 274 27086 710
rect 31226 358 31512 708
<< metal3 >>
rect 118 5146 610 5151
rect 118 4162 128 5146
rect 600 4162 610 5146
rect 118 4157 610 4162
rect 18016 3096 18262 3101
rect 18016 2740 18026 3096
rect 18252 2740 18262 3096
rect 18016 2735 18262 2740
rect 22996 2342 23316 2347
rect 17376 2321 19740 2322
rect 17376 2023 17377 2321
rect 17675 2023 19740 2321
rect 17376 2022 19740 2023
rect 20040 2022 20046 2322
rect 22996 2006 23006 2342
rect 23306 2006 23316 2342
rect 22996 2001 23316 2006
rect 26804 710 27096 715
rect 22378 670 22654 675
rect 22378 428 22388 670
rect 22644 428 22654 670
rect 22378 423 22654 428
rect 26804 274 26814 710
rect 27086 274 27096 710
rect 31216 708 31522 713
rect 31216 358 31226 708
rect 31512 358 31522 708
rect 31216 353 31522 358
rect 26804 269 27096 274
<< via3 >>
rect 128 4162 600 5146
rect 18026 2740 18252 3096
rect 17377 2023 17675 2321
rect 19740 2022 20040 2322
rect 23006 2006 23306 2342
rect 22388 428 22644 670
rect 26814 274 27086 710
rect 31226 358 31512 708
<< metal4 >>
rect 798 44952 858 45152
rect 1534 44952 1594 45152
rect 2270 44952 2330 45152
rect 3006 44952 3066 45152
rect 3742 44952 3802 45152
rect 4478 44952 4538 45152
rect 5214 44952 5274 45152
rect 5950 44952 6010 45152
rect 6686 44952 6746 45152
rect 7422 44952 7482 45152
rect 8158 44952 8218 45152
rect 8894 44952 8954 45152
rect 9630 44952 9690 45152
rect 10366 44952 10426 45152
rect 11102 44952 11162 45152
rect 11838 44952 11898 45152
rect 12574 44952 12634 45152
rect 13310 44952 13370 45152
rect 14046 44952 14106 45152
rect 14782 44952 14842 45152
rect 15518 44952 15578 45152
rect 16254 44952 16314 45152
rect 16990 44952 17050 45152
rect 17726 44952 17786 45152
rect 18462 44952 18522 45152
rect 19198 44952 19258 45152
rect 19934 44952 19994 45152
rect 20670 44952 20730 45152
rect 21406 44952 21466 45152
rect 22142 44952 22202 45152
rect 22878 44952 22938 45152
rect 23614 44952 23674 45152
rect 24350 44952 24410 45152
rect 25086 44952 25146 45152
rect 25822 44952 25882 45152
rect 26558 44952 26618 45152
rect 27294 44952 27354 45152
rect 28030 44952 28090 45152
rect 28766 44952 28826 45152
rect 29502 44952 29562 45152
rect 30238 44952 30298 45152
rect 30974 44952 31034 45152
rect 31710 44952 31770 45152
rect 200 5147 500 44152
rect 127 5146 601 5147
rect 127 4162 128 5146
rect 600 4162 601 5146
rect 127 4161 601 4162
rect 200 1000 500 4161
rect 9800 2322 10100 44152
rect 18025 3096 18253 3097
rect 18025 2740 18026 3096
rect 18252 2740 18253 3096
rect 18025 2739 18253 2740
rect 9800 2321 17676 2322
rect 9800 2023 17377 2321
rect 17675 2023 17676 2321
rect 9800 2022 17676 2023
rect 9800 1000 10100 2022
rect 400 0 520 200
rect 4816 0 4936 200
rect 9232 0 9352 200
rect 13648 0 13768 200
rect 18064 0 18184 2739
rect 23005 2342 23307 2343
rect 19739 2322 20041 2323
rect 23005 2322 23006 2342
rect 19739 2022 19740 2322
rect 20040 2022 23006 2322
rect 19739 2021 20041 2022
rect 23005 2006 23006 2022
rect 23306 2006 23307 2342
rect 23005 2005 23307 2006
rect 26813 710 27087 711
rect 22387 670 22645 671
rect 22387 428 22388 670
rect 22644 428 22645 670
rect 22387 427 22645 428
rect 22480 0 22600 427
rect 26813 274 26814 710
rect 27086 274 27087 710
rect 31225 708 31513 709
rect 31225 358 31226 708
rect 31512 358 31513 708
rect 31225 357 31513 358
rect 26813 273 27087 274
rect 26896 0 27016 273
rect 31312 0 31432 357
use pfd  pfd_0 ~/pll/magic
timestamp 1709721316
transform -1 0 26992 0 1 4272
box 656 -1968 4324 608
<< labels >>
flabel metal4 s 30974 44952 31034 45152 0 FreeSans 480 90 0 0 clk
port 0 nsew signal input
flabel metal4 s 31710 44952 31770 45152 0 FreeSans 480 90 0 0 ena
port 1 nsew signal input
flabel metal4 s 30238 44952 30298 45152 0 FreeSans 480 90 0 0 rst_n
port 2 nsew signal input
flabel metal4 s 31312 0 31432 200 0 FreeSans 960 0 0 0 ua[0]
port 3 nsew signal bidirectional
flabel metal4 s 26896 0 27016 200 0 FreeSans 960 0 0 0 ua[1]
port 4 nsew signal bidirectional
flabel metal4 s 22480 0 22600 200 0 FreeSans 960 0 0 0 ua[2]
port 5 nsew signal bidirectional
flabel metal4 s 18064 0 18184 200 0 FreeSans 960 0 0 0 ua[3]
port 6 nsew signal bidirectional
flabel metal4 s 13648 0 13768 200 0 FreeSans 960 0 0 0 ua[4]
port 7 nsew signal bidirectional
flabel metal4 s 9232 0 9352 200 0 FreeSans 960 0 0 0 ua[5]
port 8 nsew signal bidirectional
flabel metal4 s 4816 0 4936 200 0 FreeSans 960 0 0 0 ua[6]
port 9 nsew signal bidirectional
flabel metal4 s 400 0 520 200 0 FreeSans 960 0 0 0 ua[7]
port 10 nsew signal bidirectional
flabel metal4 s 29502 44952 29562 45152 0 FreeSans 480 90 0 0 ui_in[0]
port 11 nsew signal input
flabel metal4 s 28766 44952 28826 45152 0 FreeSans 480 90 0 0 ui_in[1]
port 12 nsew signal input
flabel metal4 s 28030 44952 28090 45152 0 FreeSans 480 90 0 0 ui_in[2]
port 13 nsew signal input
flabel metal4 s 27294 44952 27354 45152 0 FreeSans 480 90 0 0 ui_in[3]
port 14 nsew signal input
flabel metal4 s 26558 44952 26618 45152 0 FreeSans 480 90 0 0 ui_in[4]
port 15 nsew signal input
flabel metal4 s 25822 44952 25882 45152 0 FreeSans 480 90 0 0 ui_in[5]
port 16 nsew signal input
flabel metal4 s 25086 44952 25146 45152 0 FreeSans 480 90 0 0 ui_in[6]
port 17 nsew signal input
flabel metal4 s 24350 44952 24410 45152 0 FreeSans 480 90 0 0 ui_in[7]
port 18 nsew signal input
flabel metal4 s 23614 44952 23674 45152 0 FreeSans 480 90 0 0 uio_in[0]
port 19 nsew signal input
flabel metal4 s 22878 44952 22938 45152 0 FreeSans 480 90 0 0 uio_in[1]
port 20 nsew signal input
flabel metal4 s 22142 44952 22202 45152 0 FreeSans 480 90 0 0 uio_in[2]
port 21 nsew signal input
flabel metal4 s 21406 44952 21466 45152 0 FreeSans 480 90 0 0 uio_in[3]
port 22 nsew signal input
flabel metal4 s 20670 44952 20730 45152 0 FreeSans 480 90 0 0 uio_in[4]
port 23 nsew signal input
flabel metal4 s 19934 44952 19994 45152 0 FreeSans 480 90 0 0 uio_in[5]
port 24 nsew signal input
flabel metal4 s 19198 44952 19258 45152 0 FreeSans 480 90 0 0 uio_in[6]
port 25 nsew signal input
flabel metal4 s 18462 44952 18522 45152 0 FreeSans 480 90 0 0 uio_in[7]
port 26 nsew signal input
flabel metal4 s 5950 44952 6010 45152 0 FreeSans 480 90 0 0 uio_oe[0]
port 27 nsew signal output
flabel metal4 s 5214 44952 5274 45152 0 FreeSans 480 90 0 0 uio_oe[1]
port 28 nsew signal output
flabel metal4 s 4478 44952 4538 45152 0 FreeSans 480 90 0 0 uio_oe[2]
port 29 nsew signal output
flabel metal4 s 3742 44952 3802 45152 0 FreeSans 480 90 0 0 uio_oe[3]
port 30 nsew signal output
flabel metal4 s 3006 44952 3066 45152 0 FreeSans 480 90 0 0 uio_oe[4]
port 31 nsew signal output
flabel metal4 s 2270 44952 2330 45152 0 FreeSans 480 90 0 0 uio_oe[5]
port 32 nsew signal output
flabel metal4 s 1534 44952 1594 45152 0 FreeSans 480 90 0 0 uio_oe[6]
port 33 nsew signal output
flabel metal4 s 798 44952 858 45152 0 FreeSans 480 90 0 0 uio_oe[7]
port 34 nsew signal output
flabel metal4 s 11838 44952 11898 45152 0 FreeSans 480 90 0 0 uio_out[0]
port 35 nsew signal output
flabel metal4 s 11102 44952 11162 45152 0 FreeSans 480 90 0 0 uio_out[1]
port 36 nsew signal output
flabel metal4 s 10366 44952 10426 45152 0 FreeSans 480 90 0 0 uio_out[2]
port 37 nsew signal output
flabel metal4 s 9630 44952 9690 45152 0 FreeSans 480 90 0 0 uio_out[3]
port 38 nsew signal output
flabel metal4 s 8894 44952 8954 45152 0 FreeSans 480 90 0 0 uio_out[4]
port 39 nsew signal output
flabel metal4 s 8158 44952 8218 45152 0 FreeSans 480 90 0 0 uio_out[5]
port 40 nsew signal output
flabel metal4 s 7422 44952 7482 45152 0 FreeSans 480 90 0 0 uio_out[6]
port 41 nsew signal output
flabel metal4 s 6686 44952 6746 45152 0 FreeSans 480 90 0 0 uio_out[7]
port 42 nsew signal output
flabel metal4 s 17726 44952 17786 45152 0 FreeSans 480 90 0 0 uo_out[0]
port 43 nsew signal output
flabel metal4 s 16990 44952 17050 45152 0 FreeSans 480 90 0 0 uo_out[1]
port 44 nsew signal output
flabel metal4 s 16254 44952 16314 45152 0 FreeSans 480 90 0 0 uo_out[2]
port 45 nsew signal output
flabel metal4 s 15518 44952 15578 45152 0 FreeSans 480 90 0 0 uo_out[3]
port 46 nsew signal output
flabel metal4 s 14782 44952 14842 45152 0 FreeSans 480 90 0 0 uo_out[4]
port 47 nsew signal output
flabel metal4 s 14046 44952 14106 45152 0 FreeSans 480 90 0 0 uo_out[5]
port 48 nsew signal output
flabel metal4 s 13310 44952 13370 45152 0 FreeSans 480 90 0 0 uo_out[6]
port 49 nsew signal output
flabel metal4 s 12574 44952 12634 45152 0 FreeSans 480 90 0 0 uo_out[7]
port 50 nsew signal output
flabel metal4 200 1000 500 44152 1 FreeSans 2 0 0 0 VPWR
port 51 nsew power bidirectional
flabel metal4 9800 1000 10100 44152 1 FreeSans 2 0 0 0 VGND
port 52 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 66976 45152
<< end >>
