* NGSPICE file created from pfd.ext - technology: sky130A

.subckt sky130_fd_sc_hd__dfrbp_2 CLK D RESET_B VGND VNB VPB VPWR Q Q_N a_1462_47#
+ a_543_47# a_651_413# a_193_47# a_805_47# a_448_47# a_639_47# a_1283_21# a_761_289#
+ a_1108_47# a_1217_47# a_1659_47# a_1270_413# a_27_47#
X0 a_1217_47# a_27_47# a_1108_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X1 a_805_47# a_761_289# a_639_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X2 a_1108_47# a_193_47# a_761_289# VNB sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X3 a_1283_21# a_1108_47# a_1462_47# VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X4 Q_N a_1659_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 a_651_413# a_27_47# a_543_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X6 VGND RESET_B a_805_47# VNB sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X7 VPWR a_1283_21# Q VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.155 ps=1.31 w=1 l=0.15
X8 VPWR CLK a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X9 a_448_47# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X10 VPWR a_1283_21# a_1659_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1522 pd=1.335 as=0.1664 ps=1.8 w=0.64 l=0.15
X11 a_761_289# a_543_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X12 VGND a_1283_21# a_1659_47# VNB sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.1092 ps=1.36 w=0.42 l=0.15
X13 a_193_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X14 a_1108_47# a_27_47# a_761_289# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X15 VPWR a_1659_47# Q_N VPB sky130_fd_pr__pfet_01v8_hvt ad=0.31 pd=2.62 as=0.135 ps=1.27 w=1 l=0.15
X16 a_543_47# a_27_47# a_448_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X17 a_1462_47# RESET_B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X18 VGND a_1659_47# Q_N VNB sky130_fd_pr__nfet_01v8 ad=0.2015 pd=1.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X19 a_543_47# a_193_47# a_448_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X20 a_448_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X21 VPWR a_1283_21# a_1270_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X22 VPWR a_1108_47# a_1283_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1197 pd=1.41 as=0.0567 ps=0.69 w=0.42 l=0.15
X23 a_1270_413# a_193_47# a_1108_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X24 a_193_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X25 a_1283_21# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X26 Q a_1283_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.10025 ps=0.985 w=0.65 l=0.15
X27 VPWR a_761_289# a_651_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X28 VGND a_1283_21# Q VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10075 ps=0.96 w=0.65 l=0.15
X29 Q_N a_1659_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X30 Q a_1283_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.1522 ps=1.335 w=1 l=0.15
X31 a_639_47# a_193_47# a_543_47# VNB sky130_fd_pr__nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X32 VGND a_1283_21# a_1217_47# VNB sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X33 a_651_413# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X34 VGND CLK a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X35 a_761_289# a_543_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
C0 VGND a_27_47# 0.253971f
C1 a_193_47# a_1217_47# 2.36e-20
C2 VPB CLK 0.069345f
C3 RESET_B a_193_47# 0.026903f
C4 a_543_47# a_761_289# 0.209641f
C5 a_1659_47# a_1283_21# 0.303605f
C6 VPWR a_761_289# 0.10497f
C7 a_1659_47# VGND 0.13852f
C8 a_1108_47# a_761_289# 0.051162f
C9 a_761_289# a_639_47# 3.16e-19
C10 VGND a_1283_21# 0.2208f
C11 RESET_B VPB 0.138482f
C12 VPB a_193_47# 0.170861f
C13 a_543_47# a_805_47# 0.001705f
C14 RESET_B a_1462_47# 0.002879f
C15 VPWR Q_N 0.157089f
C16 a_27_47# a_761_289# 0.07009f
C17 a_761_289# a_651_413# 0.097745f
C18 VPWR CLK 0.017406f
C19 a_1108_47# Q_N 1.34e-19
C20 Q_N Q 0.0061f
C21 RESET_B D 4.72e-19
C22 RESET_B a_543_47# 0.153272f
C23 a_193_47# D 0.217945f
C24 a_1283_21# a_761_289# 3.17e-21
C25 a_543_47# a_193_47# 0.229804f
C26 RESET_B a_448_47# 2.45e-19
C27 a_27_47# Q_N 1.53e-20
C28 RESET_B VPWR 0.065186f
C29 a_1108_47# a_1217_47# 0.007416f
C30 VGND a_761_289# 0.073384f
C31 a_27_47# CLK 0.233602f
C32 a_193_47# a_448_47# 0.064178f
C33 RESET_B a_1108_47# 0.236601f
C34 VPWR a_193_47# 0.395736f
C35 a_1108_47# a_193_47# 0.125324f
C36 a_1659_47# Q_N 0.145144f
C37 a_1270_413# a_761_289# 2.6e-19
C38 RESET_B a_639_47# 9.54e-19
C39 RESET_B Q 8.5e-19
C40 VPB D 0.137565f
C41 a_193_47# a_639_47# 2.28e-19
C42 VPB a_543_47# 0.095793f
C43 a_193_47# Q 1.19e-19
C44 a_1283_21# Q_N 0.002658f
C45 a_27_47# a_1217_47# 2.56e-19
C46 VPB a_448_47# 0.014137f
C47 VPB VPWR 0.250676f
C48 RESET_B a_27_47# 0.296336f
C49 VGND Q_N 0.142765f
C50 RESET_B a_651_413# 0.012196f
C51 VGND CLK 0.017208f
C52 VPB a_1108_47# 0.111392f
C53 a_27_47# a_193_47# 0.906454f
C54 VGND a_805_47# 0.00579f
C55 a_193_47# a_651_413# 0.034619f
C56 RESET_B a_1659_47# 0.00263f
C57 VPB Q 0.002023f
C58 a_1659_47# a_193_47# 6.89e-19
C59 a_543_47# D 7.35e-20
C60 RESET_B a_1283_21# 0.277236f
C61 VGND a_1217_47# 9.68e-19
C62 D a_448_47# 0.155634f
C63 VPB a_27_47# 0.261873f
C64 VPWR D 0.081188f
C65 RESET_B VGND 0.28755f
C66 a_1283_21# a_193_47# 0.042424f
C67 VPB a_651_413# 0.013543f
C68 a_543_47# a_448_47# 0.049827f
C69 a_543_47# VPWR 0.100285f
C70 VGND a_193_47# 0.063057f
C71 a_543_47# a_1108_47# 7.99e-20
C72 VPWR a_448_47# 0.068142f
C73 RESET_B a_1270_413# 2.06e-19
C74 a_1659_47# VPB 0.073099f
C75 VPWR a_1108_47# 0.171084f
C76 a_1270_413# a_193_47# 1.46e-19
C77 a_805_47# a_761_289# 3.69e-19
C78 a_543_47# a_639_47# 0.013793f
C79 a_639_47# a_448_47# 4.61e-19
C80 VPB a_1283_21# 0.2414f
C81 VPWR Q 0.014118f
C82 a_27_47# D 0.132849f
C83 VPB VGND 0.013806f
C84 a_543_47# a_27_47# 0.115353f
C85 a_1462_47# a_1283_21# 0.007399f
C86 a_543_47# a_651_413# 0.057222f
C87 a_761_289# a_1217_47# 4.2e-19
C88 a_27_47# a_448_47# 0.093133f
C89 RESET_B a_761_289# 0.166114f
C90 a_1462_47# VGND 0.002121f
C91 VPWR a_27_47# 0.152295f
C92 VPWR a_651_413# 0.12856f
C93 a_27_47# a_1108_47# 0.102355f
C94 a_193_47# a_761_289# 0.186387f
C95 a_1283_21# D 2.77e-22
C96 a_1659_47# VPWR 0.205837f
C97 a_27_47# a_639_47# 0.001881f
C98 a_27_47# Q 3.03e-20
C99 VGND D 0.051614f
C100 a_1283_21# a_543_47# 3.83e-21
C101 a_1659_47# a_1108_47# 0.00277f
C102 VGND a_543_47# 0.122935f
C103 a_1283_21# a_448_47# 1.11e-21
C104 a_1283_21# VPWR 0.156931f
C105 RESET_B Q_N 2.83e-19
C106 VPB a_761_289# 0.099418f
C107 a_1659_47# Q 0.185134f
C108 VGND a_448_47# 0.0661f
C109 a_1283_21# a_1108_47# 0.245854f
C110 VGND VPWR 0.096782f
C111 RESET_B CLK 1.09e-19
C112 a_27_47# a_651_413# 9.73e-19
C113 a_193_47# Q_N 9.35e-20
C114 RESET_B a_805_47# 0.003155f
C115 VGND a_1108_47# 0.147486f
C116 CLK a_193_47# 7.94e-19
C117 a_1283_21# Q 0.053245f
C118 a_1270_413# VPWR 7.19e-19
C119 a_1659_47# a_27_47# 5.63e-20
C120 VGND a_639_47# 0.008634f
C121 VGND Q 0.114874f
C122 a_1270_413# a_1108_47# 0.006453f
C123 RESET_B a_1217_47# 6.03e-19
C124 a_1283_21# a_27_47# 0.043643f
C125 VPB Q_N 0.004225f
C126 Q_N VNB 0.025191f
C127 Q VNB 0.003804f
C128 VGND VNB 1.24553f
C129 VPWR VNB 1.02447f
C130 RESET_B VNB 0.260034f
C131 D VNB 0.159894f
C132 CLK VNB 0.195254f
C133 VPB VNB 2.19949f
C134 a_1659_47# VNB 0.21348f
C135 a_651_413# VNB 0.004694f
C136 a_448_47# VNB 0.013901f
C137 a_1108_47# VNB 0.127984f
C138 a_1283_21# VNB 0.492394f
C139 a_543_47# VNB 0.157869f
C140 a_761_289# VNB 0.120848f
C141 a_193_47# VNB 0.272482f
C142 a_27_47# VNB 0.495595f
.ends

.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X a_147_75# a_61_75#
X0 X a_61_75# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.16655 ps=1.39 w=1 l=0.15
X1 VPWR a_61_75# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.38 pd=2.76 as=0.195 ps=1.39 w=1 l=0.15
X2 VPWR B a_61_75# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.16655 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X3 VGND B a_147_75# VNB sky130_fd_pr__nfet_01v8 ad=0.1118 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X4 X a_61_75# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.1118 ps=1.04 w=0.65 l=0.15
X5 VGND a_61_75# X VNB sky130_fd_pr__nfet_01v8 ad=0.247 pd=2.06 as=0.12675 ps=1.04 w=0.65 l=0.15
X6 a_61_75# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X7 a_147_75# A a_61_75# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
C0 a_61_75# a_147_75# 0.006569f
C1 VPWR X 0.194597f
C2 VPB B 0.064248f
C3 VPB a_61_75# 0.087048f
C4 VGND a_147_75# 0.004769f
C5 B A 0.096585f
C6 a_61_75# A 0.085863f
C7 VGND VPB 0.009503f
C8 VGND A 0.015556f
C9 VPWR B 0.012524f
C10 VPWR a_61_75# 0.158516f
C11 B X 0.002798f
C12 a_61_75# X 0.149596f
C13 VGND VPWR 0.07134f
C14 VGND X 0.153129f
C15 VPB A 0.08239f
C16 a_61_75# B 0.142002f
C17 VPWR a_147_75# 6.31e-19
C18 VGND B 0.011526f
C19 a_147_75# X 5.82e-19
C20 VGND a_61_75# 0.125003f
C21 VPWR VPB 0.090199f
C22 VPB X 0.005513f
C23 VPWR A 0.040281f
C24 A X 1.84e-19
C25 VGND VNB 0.390327f
C26 X VNB 0.027496f
C27 B VNB 0.111386f
C28 A VNB 0.177011f
C29 VPWR VNB 0.349659f
C30 VPB VNB 0.604764f
C31 a_61_75# VNB 0.263837f
.ends

.subckt sky130_fd_sc_hd__inv_4 A VGND VNB VPB VPWR Y
X0 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X7 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
C0 A VGND 0.081909f
C1 VPB Y 0.015896f
C2 Y VPWR 0.361779f
C3 A Y 0.359887f
C4 Y VGND 0.262586f
C5 VPB VPWR 0.065385f
C6 A VPB 0.141975f
C7 VPB VGND 0.006668f
C8 A VPWR 0.098226f
C9 VPWR VGND 0.050092f
C10 VGND VNB 0.326816f
C11 Y VNB 0.084947f
C12 VPWR VNB 0.296394f
C13 A VNB 0.451855f
C14 VPB VNB 0.516168f
.ends

 
.subckt pfd_pex VSS VDD A QA QB B
Xx1 A VDD x4/Y VSS VSS VDD VDD QA x1/Q_N x1/a_1462_47# x1/a_543_47# x1/a_651_413#
+ x1/a_193_47# x1/a_805_47# x1/a_448_47# x1/a_639_47# x1/a_1283_21# x1/a_761_289#
+ x1/a_1108_47# x1/a_1217_47# x1/a_1659_47# x1/a_1270_413# x1/a_27_47# sky130_fd_sc_hd__dfrbp_2
Xx2 QA QB VSS VSS VDD VDD x4/A x2/a_147_75# x2/a_61_75# sky130_fd_sc_hd__and2_2
Xx3 B VDD x4/Y VSS VSS VDD VDD QB x3/Q_N x3/a_1462_47# x3/a_543_47# x3/a_651_413#
+ x3/a_193_47# x3/a_805_47# x3/a_448_47# x3/a_639_47# x3/a_1283_21# x3/a_761_289#
+ x3/a_1108_47# x3/a_1217_47# x3/a_1659_47# x3/a_1270_413# x3/a_27_47# sky130_fd_sc_hd__dfrbp_2
Xx4 x4/A VSS VSS VDD VDD x4/Y sky130_fd_sc_hd__inv_4
C0 VSS x4/A 0.064922f
C1 VDD x4/Y 1.068738f
C2 x4/Y x3/a_193_47# 0.078086f
C3 x3/a_1108_47# x1/a_1283_21# 1.76e-20
C4 x1/a_448_47# x4/Y 0.006797f
C5 x4/A x1/a_1108_47# 3.75e-19
C6 x3/a_1659_47# x1/a_1659_47# 0.001065f
C7 VDD x3/a_761_289# 1.79e-20
C8 x3/a_1108_47# QB 0.003568f
C9 x1/a_27_47# x4/Y 0.021492f
C10 x3/a_27_47# x3/Q_N -4.19e-21
C11 x1/a_193_47# x3/a_1283_21# 2.6e-20
C12 QA x1/a_761_289# 3.76e-19
C13 x3/a_1108_47# x2/a_61_75# 0.001741f
C14 VSS QA 0.079436f
C15 VDD x1/Q_N -0.002396f
C16 x3/a_448_47# x4/Y 0.006088f
C17 x3/a_1270_413# QB 4.92e-20
C18 VDD B 0.037258f
C19 QA x1/a_1108_47# 0.002062f
C20 x1/a_27_47# x1/Q_N -4.19e-21
C21 B x3/a_193_47# 0.001165f
C22 x3/a_761_289# x4/Y 0.028323f
C23 x1/a_27_47# B 2.72e-20
C24 x4/A x3/a_651_413# 3.63e-19
C25 VSS x3/a_1217_47# 5.01e-20
C26 QA x1/a_1659_47# 0.084248f
C27 x3/a_27_47# x1/a_193_47# 5.26e-19
C28 x3/Q_N QB 0.076678f
C29 VDD x3/a_1108_47# 5.48e-19
C30 x3/a_448_47# B 8.04e-20
C31 x1/Q_N x4/Y 1.8e-19
C32 VDD x1/a_651_413# 4.53e-19
C33 VSS x1/a_1462_47# 2.06e-19
C34 VSS x1/a_761_289# -0.001714f
C35 VDD x3/a_1270_413# 3.44e-21
C36 B x4/Y 0.002946f
C37 x1/a_27_47# x3/a_1108_47# 2.65e-20
C38 x4/A x3/a_1283_21# 1.74e-19
C39 VDD A 0.276941f
C40 x3/a_761_289# B 1.38e-19
C41 x1/a_805_47# VDD 1.49e-19
C42 x3/a_27_47# x1/a_543_47# 1.11e-21
C43 VSS x1/a_1108_47# 4.55e-19
C44 x1/a_27_47# A 0.003469f
C45 x3/a_1108_47# x4/Y 0.015946f
C46 x3/a_27_47# x3/a_1659_47# -2.46e-20
C47 x1/a_651_413# x4/Y 0.002005f
C48 VDD x3/Q_N -0.001965f
C49 QA x3/a_1283_21# 0.002893f
C50 VSS x1/a_1659_47# -2.85e-19
C51 x3/a_1270_413# x4/Y 1.87e-19
C52 x3/a_27_47# x4/A 0.002794f
C53 x3/a_543_47# QB 2.49e-19
C54 A x4/Y 2.55e-19
C55 x1/a_805_47# x4/Y 0.001847f
C56 VSS x3/a_651_413# 1.73e-19
C57 x3/a_1659_47# x1/a_1283_21# 1.13e-19
C58 x3/Q_N x4/Y 5.72e-19
C59 VSS x2/a_147_75# 0.001305f
C60 x3/a_1659_47# QB 0.096601f
C61 VDD x1/a_193_47# 0.016797f
C62 x1/a_193_47# x3/a_193_47# 2.81e-19
C63 x4/A x1/a_1283_21# 1.59e-19
C64 A B 0.019541f
C65 x4/A QB 0.029153f
C66 VSS x3/a_1283_21# 0.005368f
C67 x4/A x2/a_61_75# 0.0135f
C68 x3/a_543_47# VDD 0.001555f
C69 VSS x3/a_639_47# 1.05e-19
C70 x3/a_1283_21# x1/a_1108_47# 2.3e-20
C71 VDD x1/a_543_47# 0.006114f
C72 QA x1/a_1283_21# 0.025993f
C73 x1/a_193_47# x4/Y 0.013597f
C74 x1/a_27_47# x3/a_543_47# 1.37e-20
C75 QA QB 0.060347f
C76 x1/a_543_47# x3/a_193_47# 4.23e-19
C77 x3/a_1659_47# VDD -4.15e-19
C78 x1/a_1659_47# x3/a_1283_21# 9.92e-21
C79 QA x2/a_61_75# -7.04e-19
C80 x1/a_27_47# x1/a_543_47# -7.77e-20
C81 x1/a_193_47# x3/a_761_289# 8.32e-21
C82 x3/a_27_47# VSS 0.001358f
C83 x3/a_543_47# x4/Y 0.019185f
C84 VDD x4/A 0.191959f
C85 x1/a_193_47# x1/Q_N 1.39e-35
C86 x4/A x3/a_193_47# 6.35e-19
C87 x3/a_27_47# x1/a_1108_47# 2.11e-20
C88 x4/Y x1/a_543_47# 0.014551f
C89 x1/a_27_47# x4/A 0.002565f
C90 x3/a_1659_47# x4/Y 0.002286f
C91 x3/a_761_289# x1/a_543_47# 3.92e-20
C92 VSS x1/a_1283_21# 0.001115f
C93 QA VDD 0.252484f
C94 x3/a_1462_47# VSS 1.7e-19
C95 x3/a_805_47# VSS 6.63e-20
C96 VSS QB 0.070345f
C97 x3/a_543_47# B 1.13e-19
C98 x4/A x4/Y 0.056933f
C99 x1/a_193_47# x3/a_1108_47# 2.82e-20
C100 x1/a_448_47# QA 2.54e-20
C101 VSS x2/a_61_75# 0.044394f
C102 VSS x1/a_639_47# 1.17e-19
C103 x1/a_27_47# QA 5.73e-19
C104 x3/a_1659_47# x1/Q_N 2.7e-20
C105 VSS x1/a_1217_47# 5.78e-20
C106 x4/A x3/a_761_289# 0.002138f
C107 x1/a_1108_47# x2/a_61_75# 0.00156f
C108 x1/a_1659_47# x1/a_1283_21# -5.68e-32
C109 x3/a_543_47# x1/a_651_413# 1.24e-21
C110 x1/a_1659_47# QB 0.002508f
C111 QA x4/Y 0.007569f
C112 VDD x1/a_1462_47# 2.14e-20
C113 x3/a_27_47# x3/a_1283_21# -1.22e-20
C114 VDD x1/a_761_289# 0.002021f
C115 VSS VDD 1.455216f
C116 x1/a_761_289# x3/a_193_47# 1.78e-20
C117 VSS x3/a_193_47# 0.002869f
C118 QA x1/Q_N 0.066369f
C119 x1/a_27_47# x1/a_761_289# -2.48e-19
C120 x3/a_1217_47# x4/Y 9.15e-20
C121 VDD x1/a_1108_47# 0.002912f
C122 x1/a_27_47# VSS 2.8e-19
C123 x2/a_147_75# QB 0.002256f
C124 x4/A x3/a_1108_47# 4.07e-20
C125 x1/a_1108_47# x3/a_193_47# 8.83e-21
C126 VDD x1/a_1270_413# 1.52e-20
C127 x4/A x1/a_651_413# 5.44e-20
C128 x1/a_1462_47# x4/Y 3.98e-19
C129 x1/a_1283_21# x3/a_1283_21# 0.001687f
C130 VDD x1/a_1659_47# 0.003868f
C131 x1/a_761_289# x4/Y 0.011692f
C132 QB x3/a_1283_21# 0.036568f
C133 VSS x4/Y 0.55527f
C134 x3/a_1283_21# x2/a_61_75# 8.96e-19
C135 x1/a_27_47# x1/a_1659_47# -2.46e-20
C136 VSS x3/a_761_289# 8.47e-19
C137 x4/Y x1/a_1108_47# 0.005587f
C138 VDD x3/a_651_413# 4.62e-20
C139 x3/a_543_47# x1/a_193_47# 3.36e-21
C140 VSS x1/Q_N 0.00477f
C141 VDD x2/a_147_75# -1.99e-19
C142 x1/a_1659_47# x4/Y 2.33e-19
C143 x3/a_27_47# QB 6.7e-19
C144 VSS B 0.003206f
C145 VDD x3/a_1283_21# 3.46e-19
C146 x3/a_651_413# x4/Y 0.008881f
C147 x3/a_543_47# x1/a_543_47# 0.001216f
C148 x1/a_27_47# x3/a_1283_21# 4.6e-20
C149 VSS x3/a_1108_47# 0.00166f
C150 x4/A x1/a_193_47# 0.002973f
C151 x1/a_1283_21# QB 0.003617f
C152 VSS x3/a_1270_413# 3e-20
C153 x1/a_1283_21# x2/a_61_75# 8.5e-19
C154 VSS A 0.003056f
C155 x3/a_27_47# VDD 0.002308f
C156 x4/Y x3/a_1283_21# 0.007804f
C157 QB x2/a_61_75# 0.06191f
C158 x3/a_543_47# x4/A 0.001072f
C159 x3/a_27_47# x3/a_193_47# -1.84e-19
C160 VSS x1/a_805_47# 6.61e-20
C161 QA x1/a_193_47# 0.001315f
C162 x3/a_27_47# x1/a_448_47# 1.92e-21
C163 x3/a_639_47# x4/Y 0.001004f
C164 x4/A x1/a_543_47# 7.24e-19
C165 x3/a_27_47# x1/a_27_47# 7.09e-19
C166 VSS x3/Q_N 0.009158f
C167 VDD x1/a_1283_21# 0.013028f
C168 x3/a_27_47# x4/Y 0.063841f
C169 VDD QB 0.394022f
C170 QA x1/a_543_47# 2.62e-19
C171 QB x3/a_193_47# 7.35e-19
C172 VDD x2/a_61_75# 0.015492f
C173 x1/a_639_47# VDD 3.79e-19
C174 x1/a_27_47# x1/a_1283_21# -1.22e-20
C175 x3/Q_N x1/a_1659_47# 5.94e-20
C176 QA x3/a_1659_47# 4.13e-19
C177 VDD x1/a_1217_47# 2.11e-20
C178 VSS x1/a_193_47# 2.63e-19
C179 x3/a_448_47# QB 2.37e-20
C180 QA x4/A 2.26e-20
C181 x1/a_1283_21# x4/Y 0.002474f
C182 x3/a_1462_47# x4/Y 6.94e-20
C183 x3/a_27_47# B 0.009415f
C184 x1/a_193_47# x1/a_1108_47# 1.42e-32
C185 x3/a_543_47# x1/a_761_289# 4.26e-20
C186 x3/a_805_47# x4/Y 5.09e-19
C187 x4/Y QB 0.050631f
C188 x3/a_543_47# VSS 0.001259f
C189 x4/Y x2/a_61_75# 9.55e-19
C190 x1/a_639_47# x4/Y 0.003447f
C191 x3/a_761_289# QB 3.38e-19
C192 x4/Y x1/a_1217_47# 3.35e-19
C193 VDD x3/a_193_47# 0.003037f
C194 VSS x1/a_543_47# -1.78e-19
C195 x1/a_448_47# VDD 0.001274f
C196 x1/Q_N QB 7.23e-19
C197 x1/a_27_47# VDD 0.041518f
C198 x1/a_448_47# x3/a_193_47# 2.61e-20
C199 VSS x3/a_1659_47# 0.006621f
C200 x1/a_27_47# x3/a_193_47# 0.001366f
C201 VDD x3/a_448_47# 7.49e-20
C202 x1/a_761_289# x4/A 0.002468f
C203 x3/a_27_47# A 5.05e-19
C204 VDD 0 9.515211f
C205 x4/A 0 0.603123f
C206 x3/Q_N 0 0.025191f
C207 QB 0 1.514412f
C208 B 0 0.71044f
C209 x3/a_1659_47# 0 0.21348f
C210 x3/a_651_413# 0 0.004694f
C211 x3/a_448_47# 0 0.013901f
C212 x3/a_1108_47# 0 0.127984f
C213 x3/a_1283_21# 0 0.492394f
C214 x3/a_543_47# 0 0.157869f
C215 x3/a_761_289# 0 0.120848f
C216 x3/a_193_47# 0 0.272482f
C217 x3/a_27_47# 0 0.495595f
C218 x2/a_61_75# 0 0.263837f
C219 x1/Q_N 0 0.025191f
C220 QA 0 1.749791f
C221 VSS 0 1.458553f
C222 x4/Y 0 1.310204f
C223 A 0 0.706987f
C224 x1/a_1659_47# 0 0.21348f
C225 x1/a_651_413# 0 0.004694f
C226 x1/a_448_47# 0 0.013901f
C227 x1/a_1108_47# 0 0.127984f
C228 x1/a_1283_21# 0 0.492394f
C229 x1/a_543_47# 0 0.157869f
C230 x1/a_761_289# 0 0.120848f
C231 x1/a_193_47# 0 0.272482f
C232 x1/a_27_47# 0 0.495595f
.ends

