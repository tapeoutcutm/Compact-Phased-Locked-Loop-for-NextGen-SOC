MACRO NFD
  CLASS BLOCK ;
  FOREIGN NFD ;
  ORIGIN -0.210 11.670 ;
  SIZE 39.330 BY 5.960 ;
  PIN VSS
    ANTENNADIFFAREA 4.153150 ;
    PORT
      LAYER pwell ;
        RECT 1.020 -9.415 2.040 -9.410 ;
        RECT 5.370 -9.415 6.280 -9.195 ;
        RECT 7.820 -9.415 11.505 -9.185 ;
        RECT 18.620 -9.365 19.530 -9.145 ;
        RECT 21.070 -9.365 24.755 -9.135 ;
        RECT 1.020 -9.460 11.505 -9.415 ;
        RECT 15.105 -9.390 24.755 -9.365 ;
        RECT 32.040 -9.385 32.950 -9.165 ;
        RECT 34.490 -9.385 38.175 -9.155 ;
        RECT 28.525 -9.390 38.175 -9.385 ;
        RECT 15.105 -9.460 38.175 -9.390 ;
        RECT 1.020 -9.960 38.175 -9.460 ;
        RECT 1.020 -10.030 24.755 -9.960 ;
        RECT 1.020 -10.095 11.505 -10.030 ;
        RECT 15.105 -10.045 24.755 -10.030 ;
        RECT 1.020 -10.140 2.165 -10.095 ;
        RECT 1.995 -10.285 2.165 -10.140 ;
        RECT 15.245 -10.235 15.415 -10.045 ;
        RECT 28.525 -10.065 38.175 -9.960 ;
        RECT 28.665 -10.255 28.835 -10.065 ;
      LAYER li1 ;
        RECT 1.160 -10.120 1.680 -9.500 ;
        RECT 2.365 -10.115 2.695 -9.735 ;
        RECT 3.305 -10.115 3.555 -9.655 ;
        RECT 5.250 -10.115 5.620 -9.615 ;
        RECT 7.435 -10.115 7.645 -9.585 ;
        RECT 8.410 -10.115 8.580 -9.505 ;
        RECT 9.250 -10.115 9.420 -9.600 ;
        RECT 10.240 -10.115 10.570 -9.375 ;
        RECT 11.165 -10.115 11.415 -9.295 ;
        RECT 15.615 -10.065 15.945 -9.685 ;
        RECT 16.555 -10.065 16.805 -9.605 ;
        RECT 18.500 -10.065 18.870 -9.565 ;
        RECT 20.685 -10.065 20.895 -9.535 ;
        RECT 21.660 -10.065 21.830 -9.455 ;
        RECT 22.500 -10.065 22.670 -9.550 ;
        RECT 23.490 -10.065 23.820 -9.325 ;
        RECT 24.415 -10.065 24.665 -9.245 ;
        RECT 1.850 -10.120 11.510 -10.115 ;
        RECT 1.160 -10.285 11.510 -10.120 ;
        RECT 15.100 -10.235 24.760 -10.065 ;
        RECT 29.035 -10.085 29.365 -9.705 ;
        RECT 29.975 -10.085 30.225 -9.625 ;
        RECT 31.920 -10.085 32.290 -9.585 ;
        RECT 34.105 -10.085 34.315 -9.555 ;
        RECT 35.080 -10.085 35.250 -9.475 ;
        RECT 35.920 -10.085 36.090 -9.570 ;
        RECT 36.910 -10.085 37.240 -9.345 ;
        RECT 37.835 -10.085 38.085 -9.265 ;
        RECT 28.520 -10.255 38.180 -10.085 ;
        RECT 1.160 -10.310 1.990 -10.285 ;
      LAYER met1 ;
        RECT 1.850 -9.970 11.510 -9.960 ;
        RECT 15.100 -9.970 24.760 -9.910 ;
        RECT 1.850 -9.990 24.760 -9.970 ;
        RECT 28.520 -9.990 38.180 -9.930 ;
        RECT 1.850 -10.030 38.180 -9.990 ;
        RECT 1.850 -10.270 39.520 -10.030 ;
        RECT 1.850 -10.390 24.760 -10.270 ;
        RECT 1.850 -10.440 11.520 -10.390 ;
        RECT 28.520 -10.400 39.520 -10.270 ;
        RECT 28.520 -10.410 38.180 -10.400 ;
        RECT 11.120 -10.450 11.520 -10.440 ;
        RECT 38.540 -10.670 39.520 -10.400 ;
        RECT 38.540 -11.670 39.540 -10.670 ;
    END
  END VSS
  PIN f0_8
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER li1 ;
        RECT 35.410 -8.595 35.740 -7.750 ;
        RECT 35.410 -8.675 35.820 -8.595 ;
        RECT 35.585 -8.725 35.820 -8.675 ;
        RECT 35.630 -9.305 35.820 -8.725 ;
        RECT 35.575 -9.345 35.820 -9.305 ;
        RECT 35.420 -9.430 35.820 -9.345 ;
        RECT 35.420 -9.865 35.750 -9.430 ;
      LAYER met1 ;
        RECT 35.000 -6.830 36.000 -5.830 ;
        RECT 35.140 -7.000 35.900 -6.830 ;
        RECT 35.220 -8.220 35.850 -7.910 ;
        RECT 35.380 -9.530 35.760 -8.220 ;
        RECT 35.390 -9.770 35.760 -9.530 ;
      LAYER met2 ;
        RECT 35.190 -7.050 35.850 -6.540 ;
        RECT 35.250 -7.920 35.810 -7.050 ;
        RECT 35.270 -8.270 35.800 -7.920 ;
    END
  END f0_8
  PIN f0_4
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER li1 ;
        RECT 21.990 -8.575 22.320 -7.730 ;
        RECT 21.990 -8.655 22.400 -8.575 ;
        RECT 22.165 -8.705 22.400 -8.655 ;
        RECT 22.210 -9.285 22.400 -8.705 ;
        RECT 22.155 -9.325 22.400 -9.285 ;
        RECT 22.000 -9.410 22.400 -9.325 ;
        RECT 22.000 -9.845 22.330 -9.410 ;
      LAYER met1 ;
        RECT 21.610 -6.830 22.610 -5.830 ;
        RECT 21.760 -6.960 22.520 -6.830 ;
        RECT 21.810 -8.180 22.440 -7.870 ;
        RECT 21.970 -9.450 22.300 -8.180 ;
        RECT 21.970 -9.760 22.340 -9.450 ;
      LAYER met2 ;
        RECT 21.810 -7.010 22.470 -6.500 ;
        RECT 21.890 -7.820 22.360 -7.010 ;
        RECT 21.860 -8.230 22.390 -7.820 ;
    END
  END f0_4
  PIN f0_2
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER li1 ;
        RECT 8.740 -8.625 9.070 -7.780 ;
        RECT 8.740 -8.705 9.150 -8.625 ;
        RECT 8.915 -8.755 9.150 -8.705 ;
        RECT 8.960 -9.335 9.150 -8.755 ;
        RECT 8.905 -9.375 9.150 -9.335 ;
        RECT 8.750 -9.460 9.150 -9.375 ;
        RECT 8.750 -9.895 9.080 -9.460 ;
      LAYER met1 ;
        RECT 8.360 -6.840 9.360 -5.840 ;
        RECT 8.470 -6.960 9.230 -6.840 ;
        RECT 8.560 -8.290 9.190 -7.980 ;
        RECT 8.690 -9.540 9.090 -8.290 ;
        RECT 8.720 -9.800 9.090 -9.540 ;
      LAYER met2 ;
        RECT 8.520 -6.920 9.180 -6.500 ;
        RECT 8.520 -7.010 9.190 -6.920 ;
        RECT 8.540 -8.000 9.190 -7.010 ;
        RECT 8.610 -8.340 9.140 -8.000 ;
    END
  END f0_2
  PIN VDD
    ANTENNADIFFAREA 5.946950 ;
    PORT
      LAYER nwell ;
        RECT 14.910 -7.260 24.950 -7.240 ;
        RECT 14.910 -7.280 39.050 -7.260 ;
        RECT 11.520 -7.290 39.050 -7.280 ;
        RECT 1.660 -8.800 39.050 -7.290 ;
        RECT 1.660 -8.830 38.370 -8.800 ;
        RECT 1.660 -8.845 24.950 -8.830 ;
        RECT 1.660 -8.870 15.070 -8.845 ;
        RECT 28.330 -8.865 38.370 -8.830 ;
        RECT 1.660 -8.895 11.700 -8.870 ;
      LAYER li1 ;
        RECT 38.130 -7.330 38.860 -7.290 ;
        RECT 1.850 -7.565 11.510 -7.395 ;
        RECT 15.100 -7.515 24.760 -7.345 ;
        RECT 38.130 -7.360 38.890 -7.330 ;
        RECT 38.030 -7.365 38.890 -7.360 ;
        RECT 2.365 -8.065 2.695 -7.565 ;
        RECT 3.290 -8.025 3.555 -7.565 ;
        RECT 5.460 -8.365 5.630 -7.565 ;
        RECT 7.340 -8.065 7.655 -7.565 ;
        RECT 8.400 -8.575 8.570 -7.565 ;
        RECT 9.240 -8.480 9.415 -7.565 ;
        RECT 10.275 -8.705 10.490 -7.565 ;
        RECT 11.165 -8.705 11.415 -7.565 ;
        RECT 15.615 -8.015 15.945 -7.515 ;
        RECT 16.540 -7.975 16.805 -7.515 ;
        RECT 18.710 -8.315 18.880 -7.515 ;
        RECT 20.590 -8.015 20.905 -7.515 ;
        RECT 21.650 -8.525 21.820 -7.515 ;
        RECT 22.490 -8.430 22.665 -7.515 ;
        RECT 23.525 -8.655 23.740 -7.515 ;
        RECT 24.415 -8.655 24.665 -7.515 ;
        RECT 28.520 -7.535 38.890 -7.365 ;
        RECT 29.035 -8.035 29.365 -7.535 ;
        RECT 29.960 -7.995 30.225 -7.535 ;
        RECT 32.130 -8.335 32.300 -7.535 ;
        RECT 34.010 -8.035 34.325 -7.535 ;
        RECT 35.070 -8.545 35.240 -7.535 ;
        RECT 35.910 -8.450 36.085 -7.535 ;
        RECT 36.945 -8.675 37.160 -7.535 ;
        RECT 37.835 -7.570 38.890 -7.535 ;
        RECT 37.835 -8.675 38.085 -7.570 ;
        RECT 38.360 -8.620 38.890 -7.570 ;
      LAYER met1 ;
        RECT 0.210 -7.230 1.210 -5.710 ;
        RECT 0.210 -7.240 2.260 -7.230 ;
        RECT 0.210 -7.250 11.510 -7.240 ;
        RECT 15.100 -7.250 24.760 -7.190 ;
        RECT 0.210 -7.290 24.760 -7.250 ;
        RECT 28.520 -7.290 38.180 -7.210 ;
        RECT 0.210 -7.570 38.180 -7.290 ;
        RECT 0.210 -7.670 24.760 -7.570 ;
        RECT 0.210 -7.700 11.510 -7.670 ;
        RECT 28.520 -7.690 38.180 -7.570 ;
        RECT 1.850 -7.720 11.510 -7.700 ;
    END
  END VDD
  PIN clk
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER li1 ;
        RECT 1.940 -8.690 2.290 -8.575 ;
        RECT 0.570 -9.190 2.290 -8.690 ;
        RECT 1.940 -9.225 2.290 -9.190 ;
      LAYER met1 ;
        RECT 0.230 -8.660 1.230 -8.460 ;
        RECT 0.230 -9.220 1.290 -8.660 ;
        RECT 0.230 -9.460 1.230 -9.220 ;
    END
  END clk
  OBS
      LAYER li1 ;
        RECT 2.025 -8.235 2.195 -7.735 ;
        RECT 2.025 -8.405 2.690 -8.235 ;
        RECT 2.460 -9.395 2.690 -8.405 ;
        RECT 2.025 -9.565 2.690 -9.395 ;
        RECT 2.025 -9.855 2.195 -9.565 ;
        RECT 2.865 -9.855 3.050 -7.735 ;
        RECT 3.725 -8.160 3.975 -7.735 ;
        RECT 4.185 -8.010 5.290 -7.840 ;
        RECT 3.670 -8.290 3.975 -8.160 ;
        RECT 3.220 -9.485 3.500 -8.535 ;
        RECT 3.670 -9.395 3.840 -8.290 ;
        RECT 4.010 -9.075 4.250 -8.480 ;
        RECT 4.420 -8.545 4.950 -8.180 ;
        RECT 4.420 -9.245 4.590 -8.545 ;
        RECT 5.120 -8.625 5.290 -8.010 ;
        RECT 5.800 -8.065 6.050 -7.735 ;
        RECT 6.275 -8.035 7.160 -7.865 ;
        RECT 5.120 -8.715 5.630 -8.625 ;
        RECT 3.670 -9.525 3.895 -9.395 ;
        RECT 4.065 -9.465 4.590 -9.245 ;
        RECT 4.760 -8.885 5.630 -8.715 ;
        RECT 3.725 -9.665 3.895 -9.525 ;
        RECT 4.760 -9.665 4.930 -8.885 ;
        RECT 5.460 -8.955 5.630 -8.885 ;
        RECT 5.140 -9.135 5.340 -9.105 ;
        RECT 5.800 -9.135 5.970 -8.065 ;
        RECT 6.140 -8.955 6.330 -8.235 ;
        RECT 5.140 -9.435 5.970 -9.135 ;
        RECT 6.500 -9.165 6.820 -8.205 ;
        RECT 3.725 -9.835 4.060 -9.665 ;
        RECT 4.255 -9.835 4.930 -9.665 ;
        RECT 5.800 -9.665 5.970 -9.435 ;
        RECT 6.355 -9.495 6.820 -9.165 ;
        RECT 6.990 -8.875 7.160 -8.035 ;
        RECT 7.890 -8.295 8.230 -7.735 ;
        RECT 7.330 -8.670 8.230 -8.295 ;
        RECT 9.755 -8.485 10.085 -7.755 ;
        RECT 8.040 -8.875 8.230 -8.670 ;
        RECT 9.815 -8.875 10.085 -8.485 ;
        RECT 10.660 -8.705 10.995 -7.735 ;
        RECT 15.275 -8.185 15.445 -7.685 ;
        RECT 15.275 -8.355 15.940 -8.185 ;
        RECT 10.780 -8.850 10.995 -8.705 ;
        RECT 6.990 -9.205 7.870 -8.875 ;
        RECT 8.040 -9.205 8.790 -8.875 ;
        RECT 9.815 -9.205 10.610 -8.875 ;
        RECT 10.780 -8.880 11.000 -8.850 ;
        RECT 15.190 -8.880 15.540 -8.525 ;
        RECT 10.780 -9.090 15.540 -8.880 ;
        RECT 10.780 -9.100 11.000 -9.090 ;
        RECT 6.990 -9.665 7.160 -9.205 ;
        RECT 8.040 -9.375 8.240 -9.205 ;
        RECT 5.800 -9.835 6.205 -9.665 ;
        RECT 6.375 -9.835 7.160 -9.665 ;
        RECT 7.910 -9.900 8.240 -9.375 ;
        RECT 9.815 -9.585 10.015 -9.205 ;
        RECT 10.780 -9.315 10.995 -9.100 ;
        RECT 15.190 -9.175 15.540 -9.090 ;
        RECT 9.755 -9.855 10.015 -9.585 ;
        RECT 10.740 -9.935 10.995 -9.315 ;
        RECT 15.710 -9.345 15.940 -8.355 ;
        RECT 15.275 -9.515 15.940 -9.345 ;
        RECT 15.275 -9.805 15.445 -9.515 ;
        RECT 16.115 -9.805 16.300 -7.685 ;
        RECT 16.975 -8.110 17.225 -7.685 ;
        RECT 17.435 -7.960 18.540 -7.790 ;
        RECT 16.920 -8.240 17.225 -8.110 ;
        RECT 16.470 -9.435 16.750 -8.485 ;
        RECT 16.920 -9.345 17.090 -8.240 ;
        RECT 17.260 -9.025 17.500 -8.430 ;
        RECT 17.670 -8.495 18.200 -8.130 ;
        RECT 17.670 -9.195 17.840 -8.495 ;
        RECT 18.370 -8.575 18.540 -7.960 ;
        RECT 19.050 -8.015 19.300 -7.685 ;
        RECT 19.525 -7.985 20.410 -7.815 ;
        RECT 18.370 -8.665 18.880 -8.575 ;
        RECT 16.920 -9.475 17.145 -9.345 ;
        RECT 17.315 -9.415 17.840 -9.195 ;
        RECT 18.010 -8.835 18.880 -8.665 ;
        RECT 16.975 -9.615 17.145 -9.475 ;
        RECT 18.010 -9.615 18.180 -8.835 ;
        RECT 18.710 -8.905 18.880 -8.835 ;
        RECT 18.390 -9.085 18.590 -9.055 ;
        RECT 19.050 -9.085 19.220 -8.015 ;
        RECT 19.390 -8.905 19.580 -8.185 ;
        RECT 18.390 -9.385 19.220 -9.085 ;
        RECT 19.750 -9.115 20.070 -8.155 ;
        RECT 16.975 -9.785 17.310 -9.615 ;
        RECT 17.505 -9.785 18.180 -9.615 ;
        RECT 19.050 -9.615 19.220 -9.385 ;
        RECT 19.605 -9.445 20.070 -9.115 ;
        RECT 20.240 -8.825 20.410 -7.985 ;
        RECT 21.140 -8.245 21.480 -7.685 ;
        RECT 20.580 -8.620 21.480 -8.245 ;
        RECT 23.005 -8.435 23.335 -7.705 ;
        RECT 21.290 -8.825 21.480 -8.620 ;
        RECT 23.065 -8.825 23.335 -8.435 ;
        RECT 23.910 -8.655 24.245 -7.685 ;
        RECT 28.695 -8.205 28.865 -7.705 ;
        RECT 28.695 -8.375 29.360 -8.205 ;
        RECT 20.240 -9.155 21.120 -8.825 ;
        RECT 21.290 -9.155 22.040 -8.825 ;
        RECT 23.065 -9.155 23.860 -8.825 ;
        RECT 24.030 -8.850 24.245 -8.655 ;
        RECT 28.610 -8.850 28.960 -8.545 ;
        RECT 24.030 -9.060 28.960 -8.850 ;
        RECT 20.240 -9.615 20.410 -9.155 ;
        RECT 21.290 -9.325 21.490 -9.155 ;
        RECT 19.050 -9.785 19.455 -9.615 ;
        RECT 19.625 -9.785 20.410 -9.615 ;
        RECT 21.160 -9.850 21.490 -9.325 ;
        RECT 23.065 -9.535 23.265 -9.155 ;
        RECT 24.030 -9.265 24.245 -9.060 ;
        RECT 28.610 -9.195 28.960 -9.060 ;
        RECT 23.005 -9.805 23.265 -9.535 ;
        RECT 23.990 -9.885 24.245 -9.265 ;
        RECT 29.130 -9.365 29.360 -8.375 ;
        RECT 28.695 -9.535 29.360 -9.365 ;
        RECT 28.695 -9.825 28.865 -9.535 ;
        RECT 29.535 -9.825 29.720 -7.705 ;
        RECT 30.395 -8.130 30.645 -7.705 ;
        RECT 30.855 -7.980 31.960 -7.810 ;
        RECT 30.340 -8.260 30.645 -8.130 ;
        RECT 29.890 -9.455 30.170 -8.505 ;
        RECT 30.340 -9.365 30.510 -8.260 ;
        RECT 30.680 -9.045 30.920 -8.450 ;
        RECT 31.090 -8.515 31.620 -8.150 ;
        RECT 31.090 -9.215 31.260 -8.515 ;
        RECT 31.790 -8.595 31.960 -7.980 ;
        RECT 32.470 -8.035 32.720 -7.705 ;
        RECT 32.945 -8.005 33.830 -7.835 ;
        RECT 31.790 -8.685 32.300 -8.595 ;
        RECT 30.340 -9.495 30.565 -9.365 ;
        RECT 30.735 -9.435 31.260 -9.215 ;
        RECT 31.430 -8.855 32.300 -8.685 ;
        RECT 30.395 -9.635 30.565 -9.495 ;
        RECT 31.430 -9.635 31.600 -8.855 ;
        RECT 32.130 -8.925 32.300 -8.855 ;
        RECT 31.810 -9.105 32.010 -9.075 ;
        RECT 32.470 -9.105 32.640 -8.035 ;
        RECT 32.810 -8.925 33.000 -8.205 ;
        RECT 31.810 -9.405 32.640 -9.105 ;
        RECT 33.170 -9.135 33.490 -8.175 ;
        RECT 30.395 -9.805 30.730 -9.635 ;
        RECT 30.925 -9.805 31.600 -9.635 ;
        RECT 32.470 -9.635 32.640 -9.405 ;
        RECT 33.025 -9.465 33.490 -9.135 ;
        RECT 33.660 -8.845 33.830 -8.005 ;
        RECT 34.560 -8.265 34.900 -7.705 ;
        RECT 34.000 -8.640 34.900 -8.265 ;
        RECT 36.425 -8.455 36.755 -7.725 ;
        RECT 34.710 -8.845 34.900 -8.640 ;
        RECT 36.485 -8.845 36.755 -8.455 ;
        RECT 37.330 -8.675 37.665 -7.705 ;
        RECT 33.660 -9.175 34.540 -8.845 ;
        RECT 34.710 -9.175 35.460 -8.845 ;
        RECT 36.485 -9.175 37.280 -8.845 ;
        RECT 33.660 -9.635 33.830 -9.175 ;
        RECT 34.710 -9.345 34.910 -9.175 ;
        RECT 32.470 -9.805 32.875 -9.635 ;
        RECT 33.045 -9.805 33.830 -9.635 ;
        RECT 34.580 -9.870 34.910 -9.345 ;
        RECT 36.485 -9.555 36.685 -9.175 ;
        RECT 37.450 -9.285 37.665 -8.675 ;
        RECT 36.425 -9.825 36.685 -9.555 ;
        RECT 37.410 -9.905 37.665 -9.285 ;
      LAYER met1 ;
        RECT 15.670 -8.210 15.960 -8.165 ;
        RECT 17.770 -8.210 18.060 -8.165 ;
        RECT 19.340 -8.210 19.630 -8.165 ;
        RECT 2.420 -8.260 2.710 -8.215 ;
        RECT 4.520 -8.260 4.810 -8.215 ;
        RECT 6.090 -8.260 6.380 -8.215 ;
        RECT 2.420 -8.400 6.380 -8.260 ;
        RECT 15.670 -8.350 19.630 -8.210 ;
        RECT 15.670 -8.395 15.960 -8.350 ;
        RECT 17.770 -8.395 18.060 -8.350 ;
        RECT 19.340 -8.395 19.630 -8.350 ;
        RECT 29.090 -8.230 29.380 -8.185 ;
        RECT 31.190 -8.230 31.480 -8.185 ;
        RECT 32.760 -8.230 33.050 -8.185 ;
        RECT 29.090 -8.370 33.050 -8.230 ;
        RECT 2.420 -8.445 2.710 -8.400 ;
        RECT 4.520 -8.445 4.810 -8.400 ;
        RECT 6.090 -8.445 6.380 -8.400 ;
        RECT 29.090 -8.415 29.380 -8.370 ;
        RECT 31.190 -8.415 31.480 -8.370 ;
        RECT 32.760 -8.415 33.050 -8.370 ;
        RECT 16.065 -8.550 16.355 -8.505 ;
        RECT 17.255 -8.550 17.545 -8.505 ;
        RECT 19.775 -8.550 20.065 -8.505 ;
        RECT 2.815 -8.600 3.105 -8.555 ;
        RECT 4.005 -8.600 4.295 -8.555 ;
        RECT 6.525 -8.600 6.815 -8.555 ;
        RECT 2.815 -8.740 6.815 -8.600 ;
        RECT 16.065 -8.690 20.065 -8.550 ;
        RECT 16.065 -8.735 16.355 -8.690 ;
        RECT 17.255 -8.735 17.545 -8.690 ;
        RECT 19.775 -8.735 20.065 -8.690 ;
        RECT 29.485 -8.570 29.775 -8.525 ;
        RECT 30.675 -8.570 30.965 -8.525 ;
        RECT 33.195 -8.570 33.485 -8.525 ;
        RECT 29.485 -8.710 33.485 -8.570 ;
        RECT 2.815 -8.785 3.105 -8.740 ;
        RECT 4.005 -8.785 4.295 -8.740 ;
        RECT 6.525 -8.785 6.815 -8.740 ;
        RECT 10.780 -8.800 11.030 -8.790 ;
        RECT 3.430 -8.940 8.200 -8.930 ;
        RECT 3.180 -9.230 8.200 -8.940 ;
        RECT 10.430 -9.160 11.030 -8.800 ;
        RECT 16.430 -8.920 16.800 -8.870 ;
        RECT 21.000 -8.920 21.490 -8.790 ;
        RECT 16.430 -9.110 21.490 -8.920 ;
        RECT 23.680 -9.110 24.250 -8.750 ;
        RECT 29.485 -8.755 29.775 -8.710 ;
        RECT 30.675 -8.755 30.965 -8.710 ;
        RECT 33.195 -8.755 33.485 -8.710 ;
        RECT 16.430 -9.150 21.080 -9.110 ;
        RECT 24.000 -9.120 24.250 -9.110 ;
        RECT 29.850 -8.910 30.220 -8.880 ;
        RECT 34.620 -8.910 35.110 -8.860 ;
        RECT 16.430 -9.160 16.800 -9.150 ;
        RECT 29.850 -9.160 35.110 -8.910 ;
        RECT 37.140 -9.160 37.670 -8.800 ;
        RECT 29.850 -9.170 30.220 -9.160 ;
        RECT 34.620 -9.180 35.110 -9.160 ;
        RECT 37.420 -9.170 37.670 -9.160 ;
        RECT 3.430 -9.240 8.200 -9.230 ;
        RECT 7.710 -9.250 8.200 -9.240 ;
      LAYER met2 ;
        RECT 10.480 -8.810 10.760 -8.750 ;
        RECT 8.680 -8.870 9.090 -8.810 ;
        RECT 10.420 -8.870 10.760 -8.810 ;
        RECT 8.110 -8.880 10.760 -8.870 ;
        RECT 7.760 -9.200 10.760 -8.880 ;
        RECT 21.050 -8.790 21.440 -8.740 ;
        RECT 23.730 -8.790 24.010 -8.700 ;
        RECT 21.050 -9.080 24.010 -8.790 ;
        RECT 21.050 -9.160 21.440 -9.080 ;
        RECT 23.730 -9.160 24.010 -9.080 ;
        RECT 34.670 -8.840 35.060 -8.810 ;
        RECT 34.670 -8.850 36.780 -8.840 ;
        RECT 37.190 -8.850 37.470 -8.750 ;
        RECT 34.670 -9.160 37.470 -8.850 ;
        RECT 7.760 -9.250 8.200 -9.200 ;
        RECT 8.690 -9.210 10.760 -9.200 ;
        RECT 34.670 -9.170 36.780 -9.160 ;
        RECT 8.690 -9.250 9.090 -9.210 ;
        RECT 34.670 -9.230 35.060 -9.170 ;
        RECT 37.190 -9.210 37.470 -9.160 ;
        RECT 7.760 -9.300 8.150 -9.250 ;
  END
END NFD
END LIBRARY

