magic
tech sky130A
magscale 1 2
timestamp 1712816020
<< nwell >>
rect 1636 -376 1892 -162
rect 4192 -368 4494 -160
rect 6586 -260 6794 -38
<< pwell >>
rect 1640 -614 1822 -436
rect 4202 -602 4384 -424
rect 6582 -608 6764 -430
<< psubdiff >>
rect 1666 -512 1796 -462
rect 1666 -546 1713 -512
rect 1747 -546 1796 -512
rect 1666 -588 1796 -546
rect 4228 -500 4358 -450
rect 4228 -534 4275 -500
rect 4309 -534 4358 -500
rect 4228 -576 4358 -534
rect 6608 -506 6738 -456
rect 6608 -540 6655 -506
rect 6689 -540 6738 -506
rect 6608 -582 6738 -540
<< nsubdiff >>
rect 6632 -133 6712 -80
rect 6632 -167 6654 -133
rect 6688 -167 6712 -133
rect 1670 -250 1778 -200
rect 1670 -284 1699 -250
rect 1733 -284 1778 -250
rect 1670 -340 1778 -284
rect 4232 -240 4344 -200
rect 6632 -224 6712 -167
rect 4232 -274 4266 -240
rect 4300 -274 4344 -240
rect 4232 -322 4344 -274
<< psubdiffcont >>
rect 1713 -546 1747 -512
rect 4275 -534 4309 -500
rect 6655 -540 6689 -506
<< nsubdiffcont >>
rect 6654 -167 6688 -133
rect 1699 -284 1733 -250
rect 4266 -274 4300 -240
<< locali >>
rect 1568 -120 1736 -82
rect 4246 -88 4290 -86
rect 6642 -88 6696 -84
rect 1698 -208 1736 -120
rect 4136 -122 4290 -88
rect 6516 -122 6696 -88
rect 4246 -204 4290 -122
rect 6642 -133 6696 -122
rect 6642 -167 6654 -133
rect 6688 -167 6696 -133
rect 1680 -250 1766 -208
rect 1680 -284 1699 -250
rect 1733 -284 1766 -250
rect 1570 -311 1616 -306
rect 1570 -345 1576 -311
rect 1610 -345 1616 -311
rect 1680 -332 1766 -284
rect 4240 -240 4334 -204
rect 6642 -216 6696 -167
rect 4240 -274 4266 -240
rect 4300 -274 4334 -240
rect 4132 -310 4172 -308
rect 1570 -350 1616 -345
rect 4132 -344 4135 -310
rect 4169 -344 4172 -310
rect 4240 -316 4334 -274
rect 6516 -311 6554 -310
rect 4132 -346 4172 -344
rect 6516 -345 6518 -311
rect 6552 -345 6554 -311
rect 6516 -346 6554 -345
rect -90 -392 -36 -382
rect -90 -426 -80 -392
rect -46 -426 -36 -392
rect -90 -436 -36 -426
rect 174 -394 216 -390
rect 174 -428 179 -394
rect 213 -428 216 -394
rect 174 -436 216 -428
rect 2474 -391 2526 -380
rect 2474 -425 2483 -391
rect 2517 -425 2526 -391
rect 2474 -436 2526 -425
rect 2724 -401 2780 -384
rect 2724 -435 2738 -401
rect 2772 -435 2780 -401
rect 2724 -452 2780 -435
rect 4848 -395 4904 -386
rect 4848 -429 4859 -395
rect 4893 -429 4904 -395
rect 4848 -438 4904 -429
rect 5106 -395 5162 -370
rect 5106 -429 5122 -395
rect 5156 -429 5162 -395
rect 5106 -450 5162 -429
rect 1672 -512 1788 -468
rect 1278 -527 1314 -526
rect 1278 -561 1279 -527
rect 1313 -561 1314 -527
rect 1278 -562 1314 -561
rect 1672 -546 1711 -512
rect 1747 -546 1788 -512
rect 4234 -500 4350 -456
rect 1672 -584 1788 -546
rect 3836 -531 3878 -530
rect 3836 -565 3840 -531
rect 3874 -565 3878 -531
rect 3836 -566 3878 -565
rect 4234 -534 4273 -500
rect 4309 -534 4350 -500
rect 6614 -506 6730 -462
rect 6220 -530 6260 -528
rect 4234 -572 4350 -534
rect 6216 -531 6260 -530
rect 6216 -565 6221 -531
rect 6255 -565 6260 -531
rect 6216 -566 6260 -565
rect 6614 -540 6653 -506
rect 6689 -540 6730 -506
rect 6216 -568 6258 -566
rect 6614 -578 6730 -540
<< viali >>
rect 1576 -345 1610 -311
rect 4135 -344 4169 -310
rect 6518 -345 6552 -311
rect -80 -426 -46 -392
rect 179 -428 213 -394
rect 2483 -425 2517 -391
rect 2738 -435 2772 -401
rect 4859 -429 4893 -395
rect 5122 -429 5156 -395
rect 1279 -561 1313 -527
rect 1711 -546 1713 -512
rect 1713 -546 1745 -512
rect 3840 -565 3874 -531
rect 4273 -534 4275 -500
rect 4275 -534 4307 -500
rect 6221 -565 6255 -531
rect 6653 -540 6655 -506
rect 6655 -540 6687 -506
<< metal1 >>
rect -370 -154 5880 -62
rect -670 -376 -416 -256
rect 1578 -300 1612 -282
rect 1558 -311 1628 -300
rect 4130 -302 4178 -298
rect 1558 -345 1576 -311
rect 1610 -345 1628 -311
rect 1558 -356 1628 -345
rect 4120 -310 4184 -302
rect 6512 -304 6556 -282
rect 4120 -344 4135 -310
rect 4169 -340 4184 -310
rect 6504 -311 6566 -304
rect 4169 -344 4186 -340
rect 4120 -352 4186 -344
rect 6504 -345 6518 -311
rect 6552 -345 6566 -311
rect 6504 -352 6566 -345
rect -670 -392 -24 -376
rect 166 -386 238 -384
rect -670 -426 -80 -392
rect -46 -426 -24 -392
rect -670 -442 -24 -426
rect 164 -436 176 -386
rect 228 -398 238 -386
rect 1578 -388 1612 -356
rect 2468 -388 2532 -368
rect 4130 -372 4186 -352
rect 4130 -384 4916 -372
rect 1514 -389 2532 -388
rect 1514 -398 1526 -389
rect 166 -438 176 -436
rect 228 -434 1526 -398
rect 228 -438 238 -434
rect 166 -440 238 -438
rect 1514 -441 1526 -434
rect 1578 -391 2532 -389
rect 2724 -390 2800 -386
rect 1578 -425 2483 -391
rect 2517 -425 2532 -391
rect 1578 -428 2532 -425
rect 1578 -441 1612 -428
rect 1514 -442 1612 -441
rect -670 -488 -416 -442
rect 1578 -444 1612 -442
rect 2468 -448 2532 -428
rect 2720 -394 2800 -390
rect 2720 -446 2736 -394
rect 2788 -398 2800 -394
rect 3984 -393 4916 -384
rect 3984 -398 3996 -393
rect 2788 -444 3996 -398
rect 2788 -446 2800 -444
rect 2724 -454 2800 -446
rect 3984 -445 3996 -444
rect 4048 -395 4916 -393
rect 4048 -429 4859 -395
rect 4893 -429 4916 -395
rect 4048 -438 4916 -429
rect 4048 -445 4180 -438
rect 4836 -444 4916 -438
rect 5106 -395 5196 -388
rect 5106 -429 5122 -395
rect 5156 -397 5196 -395
rect 5177 -406 5196 -397
rect 6368 -402 6452 -392
rect 6512 -402 6556 -352
rect 6368 -403 6556 -402
rect 6368 -406 6384 -403
rect 3984 -454 4180 -445
rect 5106 -449 5125 -429
rect 5177 -449 6384 -406
rect 5106 -450 6384 -449
rect 5106 -458 5196 -450
rect 6368 -455 6384 -450
rect 6436 -452 6556 -403
rect 6436 -455 6452 -452
rect 6368 -466 6452 -455
rect 1260 -503 1344 -492
rect 1260 -555 1276 -503
rect 1328 -555 1344 -503
rect 1260 -561 1279 -555
rect 1313 -561 1344 -555
rect 1696 -512 1760 -502
rect 1696 -546 1711 -512
rect 1745 -546 1760 -512
rect 1696 -558 1760 -546
rect 3818 -506 3908 -494
rect 3818 -558 3837 -506
rect 3889 -558 3908 -506
rect 4258 -500 4322 -490
rect 4258 -522 4273 -500
rect 1260 -566 1344 -561
rect 1266 -568 1326 -566
rect 1698 -604 1758 -558
rect 3818 -565 3840 -558
rect 3874 -565 3908 -558
rect 3818 -570 3908 -565
rect 4246 -534 4273 -522
rect 4307 -522 4322 -500
rect 6638 -506 6702 -496
rect 6200 -513 6288 -506
rect 4307 -534 4330 -522
rect 3824 -572 3890 -570
rect 4246 -604 4330 -534
rect 6200 -565 6218 -513
rect 6270 -565 6288 -513
rect 6638 -532 6653 -506
rect 6200 -572 6288 -565
rect 6632 -540 6653 -532
rect 6687 -532 6702 -506
rect 6687 -540 6708 -532
rect 6204 -574 6270 -572
rect 1446 -696 5018 -604
rect 6632 -626 6708 -540
rect 6496 -672 6708 -626
rect 6632 -680 6708 -672
rect 3914 -728 4026 -726
rect 3812 -740 4112 -728
rect 1246 -765 1358 -760
rect 1246 -817 1276 -765
rect 1328 -768 1358 -765
rect 1444 -768 1544 -748
rect 1328 -816 1544 -768
rect 3812 -792 3839 -740
rect 3891 -792 4112 -740
rect 6376 -752 6486 -736
rect 3812 -804 4112 -792
rect 3998 -816 4112 -804
rect 6188 -761 6486 -752
rect 6188 -813 6219 -761
rect 6271 -813 6486 -761
rect 1328 -817 1358 -816
rect 1246 -822 1358 -817
rect 1444 -830 1544 -816
rect 6188 -820 6486 -813
rect 6188 -822 6400 -820
<< via1 >>
rect 176 -394 228 -386
rect 176 -428 179 -394
rect 179 -428 213 -394
rect 213 -428 228 -394
rect 176 -438 228 -428
rect 1526 -441 1578 -389
rect 2736 -401 2788 -394
rect 2736 -435 2738 -401
rect 2738 -435 2772 -401
rect 2772 -435 2788 -401
rect 2736 -446 2788 -435
rect 3996 -445 4048 -393
rect 5125 -429 5156 -397
rect 5156 -429 5177 -397
rect 5125 -449 5177 -429
rect 6384 -455 6436 -403
rect 1276 -527 1328 -503
rect 1276 -555 1279 -527
rect 1279 -555 1313 -527
rect 1313 -555 1328 -527
rect 3837 -531 3889 -506
rect 3837 -558 3840 -531
rect 3840 -558 3874 -531
rect 3874 -558 3889 -531
rect 6218 -531 6270 -513
rect 6218 -565 6221 -531
rect 6221 -565 6255 -531
rect 6255 -565 6270 -531
rect 1276 -817 1328 -765
rect 3839 -792 3891 -740
rect 6219 -813 6271 -761
<< metal2 >>
rect 176 -386 228 -374
rect 176 -450 228 -438
rect 1524 -389 1580 -378
rect 1524 -441 1526 -389
rect 1578 -441 1580 -389
rect 1524 -452 1580 -441
rect 2734 -394 2790 -376
rect 2734 -446 2736 -394
rect 2788 -446 2790 -394
rect 2734 -464 2790 -446
rect 3994 -393 4050 -374
rect 3994 -445 3996 -393
rect 4048 -445 4050 -393
rect 3994 -464 4050 -445
rect 5116 -397 5186 -378
rect 5116 -449 5125 -397
rect 5177 -449 5186 -397
rect 5116 -468 5186 -449
rect 6378 -403 6442 -382
rect 6378 -455 6384 -403
rect 6436 -455 6442 -403
rect 6378 -476 6442 -455
rect 1270 -503 1334 -482
rect 1270 -546 1276 -503
rect 1268 -555 1276 -546
rect 1328 -555 1334 -503
rect 1268 -576 1334 -555
rect 3828 -506 3898 -484
rect 3828 -558 3837 -506
rect 3889 -558 3898 -506
rect 3828 -574 3898 -558
rect 6210 -513 6278 -496
rect 6210 -565 6218 -513
rect 6270 -565 6278 -513
rect 1268 -750 1332 -576
rect 3828 -718 3900 -574
rect 6210 -576 6278 -565
rect 3822 -740 3908 -718
rect 1256 -765 1348 -750
rect 1256 -817 1276 -765
rect 1328 -817 1348 -765
rect 3822 -792 3839 -740
rect 3891 -792 3908 -740
rect 6208 -742 6278 -576
rect 3822 -814 3908 -792
rect 6198 -761 6292 -742
rect 6198 -813 6219 -761
rect 6271 -813 6292 -761
rect 1256 -832 1348 -817
rect 6198 -832 6292 -813
use sky130_fd_sc_hd__dfxbp_1  x1
timestamp 1712816020
transform 1 0 -110 0 1 -648
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxbp_1  x2
timestamp 1712816020
transform 1 0 2450 0 1 -650
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxbp_1  x3
timestamp 1712816020
transform 1 0 4832 0 1 -650
box -38 -48 1786 592
<< labels >>
flabel metal1 s -370 -154 5880 -62 0 FreeSans 782 0 0 0 VDD
port 1 nsew
flabel metal1 s 1446 -696 5018 -604 0 FreeSans 782 0 0 0 VSS
port 2 nsew
flabel metal1 s -670 -488 -416 -256 0 FreeSans 782 0 0 0 f0
port 3 nsew
flabel metal1 s 1444 -830 1544 -748 0 FreeSans 782 0 0 0 f0_2
port 4 nsew
flabel metal1 s 3998 -816 4112 -728 0 FreeSans 782 0 0 0 f0_4
port 5 nsew
flabel metal1 s 6376 -820 6486 -736 0 FreeSans 782 0 0 0 f0_8
port 6 nsew
<< end >>
